`include "controlFSM.sv"
`include "datapath.sv"
`include "memory.sv"

module fc_16_8_16_1_16(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 16;
	parameter N = 8;
	parameter T = 16;
	parameter R = 1;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned [3 : 0] sel;

	logic signed [T-1 : 0] parallel_out0;
	logic signed [T-1 : 0] parallel_out1;
	logic signed [T-1 : 0] parallel_out2;
	logic signed [T-1 : 0] parallel_out3;
	logic signed [T-1 : 0] parallel_out4;
	logic signed [T-1 : 0] parallel_out5;
	logic signed [T-1 : 0] parallel_out6;
	logic signed [T-1 : 0] parallel_out7;
	logic signed [T-1 : 0] parallel_out8;
	logic signed [T-1 : 0] parallel_out9;
	logic signed [T-1 : 0] parallel_out10;
	logic signed [T-1 : 0] parallel_out11;
	logic signed [T-1 : 0] parallel_out12;
	logic signed [T-1 : 0] parallel_out13;
	logic signed [T-1 : 0] parallel_out14;
	logic signed [T-1 : 0] parallel_out15;

	logic unsigned[2 : 0] addr_x;
	logic signed [15 : 0] v_out;
	logic unsigned wr_en_x;

	logic unsigned[6 : 0] addr;

	logic unsigned[6 : 0] addr_w0;
	logic signed [15 : 0] m_out0;

	logic unsigned[6 : 0] addr_w1;
	logic signed [15 : 0] m_out1;

	logic unsigned[6 : 0] addr_w2;
	logic signed [15 : 0] m_out2;

	logic unsigned[6 : 0] addr_w3;
	logic signed [15 : 0] m_out3;

	logic unsigned[6 : 0] addr_w4;
	logic signed [15 : 0] m_out4;

	logic unsigned[6 : 0] addr_w5;
	logic signed [15 : 0] m_out5;

	logic unsigned[6 : 0] addr_w6;
	logic signed [15 : 0] m_out6;

	logic unsigned[6 : 0] addr_w7;
	logic signed [15 : 0] m_out7;

	logic unsigned[6 : 0] addr_w8;
	logic signed [15 : 0] m_out8;

	logic unsigned[6 : 0] addr_w9;
	logic signed [15 : 0] m_out9;

	logic unsigned[6 : 0] addr_w10;
	logic signed [15 : 0] m_out10;

	logic unsigned[6 : 0] addr_w11;
	logic signed [15 : 0] m_out11;

	logic unsigned[6 : 0] addr_w12;
	logic signed [15 : 0] m_out12;

	logic unsigned[6 : 0] addr_w13;
	logic signed [15 : 0] m_out13;

	logic unsigned[6 : 0] addr_w14;
	logic signed [15 : 0] m_out14;

	logic unsigned[6 : 0] addr_w15;
	logic signed [15 : 0] m_out15;

	logic unsigned clear_acc;
	logic unsigned en_acc;

	always_comb begin
		addr_w0 = addr + 0;
		addr_w1 = addr + 8;
		addr_w2 = addr + 16;
		addr_w3 = addr + 24;
		addr_w4 = addr + 32;
		addr_w5 = addr + 40;
		addr_w6 = addr + 48;
		addr_w7 = addr + 56;
		addr_w8 = addr + 64;
		addr_w9 = addr + 72;
		addr_w10 = addr + 80;
		addr_w11 = addr + 88;
		addr_w12 = addr + 96;
		addr_w13 = addr + 104;
		addr_w14 = addr + 112;
		addr_w15 = addr + 120;
	end

	controlFSM #(16,8,16) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid), .countToP(sel));

	memory #(16, 8 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	mux #(16, 16) muxMod(.parallel_out0(parallel_out0), .parallel_out1(parallel_out1), .parallel_out2(parallel_out2), .parallel_out3(parallel_out3), .parallel_out4(parallel_out4), .parallel_out5(parallel_out5), .parallel_out6(parallel_out6), .parallel_out7(parallel_out7), .parallel_out8(parallel_out8), .parallel_out9(parallel_out9), .parallel_out10(parallel_out10), .parallel_out11(parallel_out11), .parallel_out12(parallel_out12), .parallel_out13(parallel_out13), .parallel_out14(parallel_out14), .parallel_out15(parallel_out15), .sel(sel), .f(output_data));

	datapath #(16, 1) datapathMod0(.clk(clk), .reset(reset), .m_out(m_out0), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out0), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod1(.clk(clk), .reset(reset), .m_out(m_out1), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out1), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod2(.clk(clk), .reset(reset), .m_out(m_out2), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out2), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod3(.clk(clk), .reset(reset), .m_out(m_out3), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out3), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod4(.clk(clk), .reset(reset), .m_out(m_out4), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out4), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod5(.clk(clk), .reset(reset), .m_out(m_out5), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out5), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod6(.clk(clk), .reset(reset), .m_out(m_out6), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out6), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod7(.clk(clk), .reset(reset), .m_out(m_out7), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out7), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod8(.clk(clk), .reset(reset), .m_out(m_out8), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out8), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod9(.clk(clk), .reset(reset), .m_out(m_out9), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out9), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod10(.clk(clk), .reset(reset), .m_out(m_out10), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out10), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod11(.clk(clk), .reset(reset), .m_out(m_out11), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out11), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod12(.clk(clk), .reset(reset), .m_out(m_out12), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out12), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod13(.clk(clk), .reset(reset), .m_out(m_out13), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out13), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod14(.clk(clk), .reset(reset), .m_out(m_out14), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out14), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod15(.clk(clk), .reset(reset), .m_out(m_out15), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out15), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	fc_16_8_16_1_16_W_rom  matrixRom(.clk(clk),.addr0(addr_w0), .addr1(addr_w1), .addr2(addr_w2), .addr3(addr_w3), .addr4(addr_w4), .addr5(addr_w5), .addr6(addr_w6), .addr7(addr_w7), .addr8(addr_w8), .addr9(addr_w9), .addr10(addr_w10), .addr11(addr_w11), .addr12(addr_w12), .addr13(addr_w13), .addr14(addr_w14), .addr15(addr_w15), .z0(m_out0), .z1(m_out1), .z2(m_out2), .z3(m_out3), .z4(m_out4), .z5(m_out5), .z6(m_out6), .z7(m_out7), .z8(m_out8), .z9(m_out9), .z10(m_out10), .z11(m_out11), .z12(m_out12), .z13(m_out13), .z14(m_out14), .z15(m_out15));

endmodule

module mux(parallel_out0, parallel_out1, parallel_out2, parallel_out3, parallel_out4, parallel_out5, parallel_out6, parallel_out7, parallel_out8, parallel_out9, parallel_out10, parallel_out11, parallel_out12, parallel_out13, parallel_out14, parallel_out15, sel, f);
	parameter T = 16;
	parameter P = 16;

	output signed [T-1 : 0] f;
	input logic unsigned [3 : 0] sel;
	input signed [T-1 : 0] parallel_out0;
	input signed [T-1 : 0] parallel_out1;
	input signed [T-1 : 0] parallel_out2;
	input signed [T-1 : 0] parallel_out3;
	input signed [T-1 : 0] parallel_out4;
	input signed [T-1 : 0] parallel_out5;
	input signed [T-1 : 0] parallel_out6;
	input signed [T-1 : 0] parallel_out7;
	input signed [T-1 : 0] parallel_out8;
	input signed [T-1 : 0] parallel_out9;
	input signed [T-1 : 0] parallel_out10;
	input signed [T-1 : 0] parallel_out11;
	input signed [T-1 : 0] parallel_out12;
	input signed [T-1 : 0] parallel_out13;
	input signed [T-1 : 0] parallel_out14;
	input signed [T-1 : 0] parallel_out15;
	logic unsigned [P*T-1 : 0] array;
	assign  array = {parallel_out0[15 : 0], parallel_out1[15 : 0], parallel_out2[15 : 0], parallel_out3[15 : 0], parallel_out4[15 : 0], parallel_out5[15 : 0], parallel_out6[15 : 0], parallel_out7[15 : 0], parallel_out8[15 : 0], parallel_out9[15 : 0], parallel_out10[15 : 0], parallel_out11[15 : 0], parallel_out12[15 : 0], parallel_out13[15 : 0], parallel_out14[15 : 0], parallel_out15[15: 0]};

	assign f = (sel == 0) ? parallel_out0 : 
			(sel == 1) ? parallel_out1 : 
			(sel == 2) ? parallel_out2 : 
			(sel == 3) ? parallel_out3 : 
			(sel == 4) ? parallel_out4 : 
			(sel == 5) ? parallel_out5 : 
			(sel == 6) ? parallel_out6 : 
			(sel == 7) ? parallel_out7 : 
			(sel == 8) ? parallel_out8 : 
			(sel == 9) ? parallel_out9 : 
			(sel == 10) ? parallel_out10 : 
			(sel == 11) ? parallel_out11 : 
			(sel == 12) ? parallel_out12 : 
			(sel == 13) ? parallel_out13 : 
			(sel == 14) ? parallel_out14 : 
			(sel == 15) ? parallel_out15 : 16'bz;
endmodule

module fc_16_8_16_1_16_W_rom(clk, addr0, addr1, addr2, addr3, addr4, addr5, addr6, addr7, addr8, addr9, addr10, addr11, addr12, addr13, addr14, addr15, z0, z1, z2, z3, z4, z5, z6, z7, z8, z9, z10, z11, z12, z13, z14, z15);
	input clk;
	input [6:0] addr0;
	input [6:0] addr1;
	input [6:0] addr2;
	input [6:0] addr3;
	input [6:0] addr4;
	input [6:0] addr5;
	input [6:0] addr6;
	input [6:0] addr7;
	input [6:0] addr8;
	input [6:0] addr9;
	input [6:0] addr10;
	input [6:0] addr11;
	input [6:0] addr12;
	input [6:0] addr13;
	input [6:0] addr14;
	input [6:0] addr15;
	output logic signed [15:0] z0;
	output logic signed [15:0] z1;
	output logic signed [15:0] z2;
	output logic signed [15:0] z3;
	output logic signed [15:0] z4;
	output logic signed [15:0] z5;
	output logic signed [15:0] z6;
	output logic signed [15:0] z7;
	output logic signed [15:0] z8;
	output logic signed [15:0] z9;
	output logic signed [15:0] z10;
	output logic signed [15:0] z11;
	output logic signed [15:0] z12;
	output logic signed [15:0] z13;
	output logic signed [15:0] z14;
	output logic signed [15:0] z15;
	always_ff @(posedge clk) begin
		case(addr0)
		0: z0 <= 16'd74;
		1: z0 <= 16'd120;
		2: z0 <= 16'd39;
		3: z0 <= -16'd125;
		4: z0 <= 16'd69;
		5: z0 <= -16'd26;
		6: z0 <= -16'd115;
		7: z0 <= -16'd84;
		8: z0 <= -16'd123;
		9: z0 <= 16'd107;
		10: z0 <= -16'd27;
		11: z0 <= 16'd118;
		12: z0 <= 16'd88;
		13: z0 <= 16'd91;
		14: z0 <= 16'd23;
		15: z0 <= 16'd64;
		16: z0 <= -16'd103;
		17: z0 <= 16'd74;
		18: z0 <= -16'd23;
		19: z0 <= -16'd14;
		20: z0 <= -16'd60;
		21: z0 <= -16'd30;
		22: z0 <= -16'd23;
		23: z0 <= -16'd101;
		24: z0 <= 16'd14;
		25: z0 <= -16'd83;
		26: z0 <= -16'd38;
		27: z0 <= 16'd74;
		28: z0 <= -16'd90;
		29: z0 <= -16'd73;
		30: z0 <= 16'd62;
		31: z0 <= 16'd112;
		32: z0 <= -16'd81;
		33: z0 <= -16'd27;
		34: z0 <= 16'd115;
		35: z0 <= 16'd116;
		36: z0 <= 16'd76;
		37: z0 <= -16'd127;
		38: z0 <= -16'd96;
		39: z0 <= 16'd81;
		40: z0 <= 16'd108;
		41: z0 <= 16'd5;
		42: z0 <= 16'd71;
		43: z0 <= 16'd68;
		44: z0 <= -16'd32;
		45: z0 <= -16'd34;
		46: z0 <= 16'd4;
		47: z0 <= -16'd6;
		48: z0 <= -16'd87;
		49: z0 <= 16'd109;
		50: z0 <= 16'd108;
		51: z0 <= -16'd19;
		52: z0 <= -16'd49;
		53: z0 <= -16'd42;
		54: z0 <= 16'd8;
		55: z0 <= 16'd93;
		56: z0 <= 16'd3;
		57: z0 <= 16'd98;
		58: z0 <= 16'd40;
		59: z0 <= 16'd41;
		60: z0 <= -16'd103;
		61: z0 <= -16'd26;
		62: z0 <= 16'd25;
		63: z0 <= -16'd56;
		64: z0 <= 16'd75;
		65: z0 <= 16'd12;
		66: z0 <= -16'd68;
		67: z0 <= 16'd23;
		68: z0 <= 16'd13;
		69: z0 <= -16'd36;
		70: z0 <= -16'd24;
		71: z0 <= -16'd6;
		72: z0 <= 16'd98;
		73: z0 <= -16'd81;
		74: z0 <= -16'd66;
		75: z0 <= -16'd62;
		76: z0 <= 16'd14;
		77: z0 <= 16'd67;
		78: z0 <= 16'd60;
		79: z0 <= 16'd55;
		80: z0 <= 16'd48;
		81: z0 <= 16'd41;
		82: z0 <= -16'd92;
		83: z0 <= -16'd128;
		84: z0 <= 16'd127;
		85: z0 <= 16'd45;
		86: z0 <= 16'd93;
		87: z0 <= 16'd2;
		88: z0 <= 16'd15;
		89: z0 <= 16'd5;
		90: z0 <= -16'd85;
		91: z0 <= 16'd41;
		92: z0 <= 16'd107;
		93: z0 <= 16'd68;
		94: z0 <= 16'd113;
		95: z0 <= 16'd55;
		96: z0 <= -16'd48;
		97: z0 <= -16'd82;
		98: z0 <= -16'd50;
		99: z0 <= 16'd94;
		100: z0 <= 16'd10;
		101: z0 <= 16'd55;
		102: z0 <= -16'd40;
		103: z0 <= -16'd20;
		104: z0 <= 16'd102;
		105: z0 <= 16'd22;
		106: z0 <= 16'd47;
		107: z0 <= -16'd12;
		108: z0 <= -16'd39;
		109: z0 <= -16'd21;
		110: z0 <= -16'd85;
		111: z0 <= -16'd118;
		112: z0 <= -16'd108;
		113: z0 <= -16'd48;
		114: z0 <= -16'd118;
		115: z0 <= -16'd109;
		116: z0 <= 16'd125;
		117: z0 <= 16'd103;
		118: z0 <= 16'd21;
		119: z0 <= 16'd12;
		120: z0 <= -16'd19;
		121: z0 <= 16'd64;
		122: z0 <= -16'd75;
		123: z0 <= -16'd40;
		124: z0 <= 16'd4;
		125: z0 <= -16'd89;
		126: z0 <= -16'd113;
		127: z0 <= 16'd85;
		endcase
		case(addr1)
		0: z1 <= 16'd74;
		1: z1 <= 16'd120;
		2: z1 <= 16'd39;
		3: z1 <= -16'd125;
		4: z1 <= 16'd69;
		5: z1 <= -16'd26;
		6: z1 <= -16'd115;
		7: z1 <= -16'd84;
		8: z1 <= -16'd123;
		9: z1 <= 16'd107;
		10: z1 <= -16'd27;
		11: z1 <= 16'd118;
		12: z1 <= 16'd88;
		13: z1 <= 16'd91;
		14: z1 <= 16'd23;
		15: z1 <= 16'd64;
		16: z1 <= -16'd103;
		17: z1 <= 16'd74;
		18: z1 <= -16'd23;
		19: z1 <= -16'd14;
		20: z1 <= -16'd60;
		21: z1 <= -16'd30;
		22: z1 <= -16'd23;
		23: z1 <= -16'd101;
		24: z1 <= 16'd14;
		25: z1 <= -16'd83;
		26: z1 <= -16'd38;
		27: z1 <= 16'd74;
		28: z1 <= -16'd90;
		29: z1 <= -16'd73;
		30: z1 <= 16'd62;
		31: z1 <= 16'd112;
		32: z1 <= -16'd81;
		33: z1 <= -16'd27;
		34: z1 <= 16'd115;
		35: z1 <= 16'd116;
		36: z1 <= 16'd76;
		37: z1 <= -16'd127;
		38: z1 <= -16'd96;
		39: z1 <= 16'd81;
		40: z1 <= 16'd108;
		41: z1 <= 16'd5;
		42: z1 <= 16'd71;
		43: z1 <= 16'd68;
		44: z1 <= -16'd32;
		45: z1 <= -16'd34;
		46: z1 <= 16'd4;
		47: z1 <= -16'd6;
		48: z1 <= -16'd87;
		49: z1 <= 16'd109;
		50: z1 <= 16'd108;
		51: z1 <= -16'd19;
		52: z1 <= -16'd49;
		53: z1 <= -16'd42;
		54: z1 <= 16'd8;
		55: z1 <= 16'd93;
		56: z1 <= 16'd3;
		57: z1 <= 16'd98;
		58: z1 <= 16'd40;
		59: z1 <= 16'd41;
		60: z1 <= -16'd103;
		61: z1 <= -16'd26;
		62: z1 <= 16'd25;
		63: z1 <= -16'd56;
		64: z1 <= 16'd75;
		65: z1 <= 16'd12;
		66: z1 <= -16'd68;
		67: z1 <= 16'd23;
		68: z1 <= 16'd13;
		69: z1 <= -16'd36;
		70: z1 <= -16'd24;
		71: z1 <= -16'd6;
		72: z1 <= 16'd98;
		73: z1 <= -16'd81;
		74: z1 <= -16'd66;
		75: z1 <= -16'd62;
		76: z1 <= 16'd14;
		77: z1 <= 16'd67;
		78: z1 <= 16'd60;
		79: z1 <= 16'd55;
		80: z1 <= 16'd48;
		81: z1 <= 16'd41;
		82: z1 <= -16'd92;
		83: z1 <= -16'd128;
		84: z1 <= 16'd127;
		85: z1 <= 16'd45;
		86: z1 <= 16'd93;
		87: z1 <= 16'd2;
		88: z1 <= 16'd15;
		89: z1 <= 16'd5;
		90: z1 <= -16'd85;
		91: z1 <= 16'd41;
		92: z1 <= 16'd107;
		93: z1 <= 16'd68;
		94: z1 <= 16'd113;
		95: z1 <= 16'd55;
		96: z1 <= -16'd48;
		97: z1 <= -16'd82;
		98: z1 <= -16'd50;
		99: z1 <= 16'd94;
		100: z1 <= 16'd10;
		101: z1 <= 16'd55;
		102: z1 <= -16'd40;
		103: z1 <= -16'd20;
		104: z1 <= 16'd102;
		105: z1 <= 16'd22;
		106: z1 <= 16'd47;
		107: z1 <= -16'd12;
		108: z1 <= -16'd39;
		109: z1 <= -16'd21;
		110: z1 <= -16'd85;
		111: z1 <= -16'd118;
		112: z1 <= -16'd108;
		113: z1 <= -16'd48;
		114: z1 <= -16'd118;
		115: z1 <= -16'd109;
		116: z1 <= 16'd125;
		117: z1 <= 16'd103;
		118: z1 <= 16'd21;
		119: z1 <= 16'd12;
		120: z1 <= -16'd19;
		121: z1 <= 16'd64;
		122: z1 <= -16'd75;
		123: z1 <= -16'd40;
		124: z1 <= 16'd4;
		125: z1 <= -16'd89;
		126: z1 <= -16'd113;
		127: z1 <= 16'd85;
		endcase
		case(addr2)
		0: z2 <= 16'd74;
		1: z2 <= 16'd120;
		2: z2 <= 16'd39;
		3: z2 <= -16'd125;
		4: z2 <= 16'd69;
		5: z2 <= -16'd26;
		6: z2 <= -16'd115;
		7: z2 <= -16'd84;
		8: z2 <= -16'd123;
		9: z2 <= 16'd107;
		10: z2 <= -16'd27;
		11: z2 <= 16'd118;
		12: z2 <= 16'd88;
		13: z2 <= 16'd91;
		14: z2 <= 16'd23;
		15: z2 <= 16'd64;
		16: z2 <= -16'd103;
		17: z2 <= 16'd74;
		18: z2 <= -16'd23;
		19: z2 <= -16'd14;
		20: z2 <= -16'd60;
		21: z2 <= -16'd30;
		22: z2 <= -16'd23;
		23: z2 <= -16'd101;
		24: z2 <= 16'd14;
		25: z2 <= -16'd83;
		26: z2 <= -16'd38;
		27: z2 <= 16'd74;
		28: z2 <= -16'd90;
		29: z2 <= -16'd73;
		30: z2 <= 16'd62;
		31: z2 <= 16'd112;
		32: z2 <= -16'd81;
		33: z2 <= -16'd27;
		34: z2 <= 16'd115;
		35: z2 <= 16'd116;
		36: z2 <= 16'd76;
		37: z2 <= -16'd127;
		38: z2 <= -16'd96;
		39: z2 <= 16'd81;
		40: z2 <= 16'd108;
		41: z2 <= 16'd5;
		42: z2 <= 16'd71;
		43: z2 <= 16'd68;
		44: z2 <= -16'd32;
		45: z2 <= -16'd34;
		46: z2 <= 16'd4;
		47: z2 <= -16'd6;
		48: z2 <= -16'd87;
		49: z2 <= 16'd109;
		50: z2 <= 16'd108;
		51: z2 <= -16'd19;
		52: z2 <= -16'd49;
		53: z2 <= -16'd42;
		54: z2 <= 16'd8;
		55: z2 <= 16'd93;
		56: z2 <= 16'd3;
		57: z2 <= 16'd98;
		58: z2 <= 16'd40;
		59: z2 <= 16'd41;
		60: z2 <= -16'd103;
		61: z2 <= -16'd26;
		62: z2 <= 16'd25;
		63: z2 <= -16'd56;
		64: z2 <= 16'd75;
		65: z2 <= 16'd12;
		66: z2 <= -16'd68;
		67: z2 <= 16'd23;
		68: z2 <= 16'd13;
		69: z2 <= -16'd36;
		70: z2 <= -16'd24;
		71: z2 <= -16'd6;
		72: z2 <= 16'd98;
		73: z2 <= -16'd81;
		74: z2 <= -16'd66;
		75: z2 <= -16'd62;
		76: z2 <= 16'd14;
		77: z2 <= 16'd67;
		78: z2 <= 16'd60;
		79: z2 <= 16'd55;
		80: z2 <= 16'd48;
		81: z2 <= 16'd41;
		82: z2 <= -16'd92;
		83: z2 <= -16'd128;
		84: z2 <= 16'd127;
		85: z2 <= 16'd45;
		86: z2 <= 16'd93;
		87: z2 <= 16'd2;
		88: z2 <= 16'd15;
		89: z2 <= 16'd5;
		90: z2 <= -16'd85;
		91: z2 <= 16'd41;
		92: z2 <= 16'd107;
		93: z2 <= 16'd68;
		94: z2 <= 16'd113;
		95: z2 <= 16'd55;
		96: z2 <= -16'd48;
		97: z2 <= -16'd82;
		98: z2 <= -16'd50;
		99: z2 <= 16'd94;
		100: z2 <= 16'd10;
		101: z2 <= 16'd55;
		102: z2 <= -16'd40;
		103: z2 <= -16'd20;
		104: z2 <= 16'd102;
		105: z2 <= 16'd22;
		106: z2 <= 16'd47;
		107: z2 <= -16'd12;
		108: z2 <= -16'd39;
		109: z2 <= -16'd21;
		110: z2 <= -16'd85;
		111: z2 <= -16'd118;
		112: z2 <= -16'd108;
		113: z2 <= -16'd48;
		114: z2 <= -16'd118;
		115: z2 <= -16'd109;
		116: z2 <= 16'd125;
		117: z2 <= 16'd103;
		118: z2 <= 16'd21;
		119: z2 <= 16'd12;
		120: z2 <= -16'd19;
		121: z2 <= 16'd64;
		122: z2 <= -16'd75;
		123: z2 <= -16'd40;
		124: z2 <= 16'd4;
		125: z2 <= -16'd89;
		126: z2 <= -16'd113;
		127: z2 <= 16'd85;
		endcase
		case(addr3)
		0: z3 <= 16'd74;
		1: z3 <= 16'd120;
		2: z3 <= 16'd39;
		3: z3 <= -16'd125;
		4: z3 <= 16'd69;
		5: z3 <= -16'd26;
		6: z3 <= -16'd115;
		7: z3 <= -16'd84;
		8: z3 <= -16'd123;
		9: z3 <= 16'd107;
		10: z3 <= -16'd27;
		11: z3 <= 16'd118;
		12: z3 <= 16'd88;
		13: z3 <= 16'd91;
		14: z3 <= 16'd23;
		15: z3 <= 16'd64;
		16: z3 <= -16'd103;
		17: z3 <= 16'd74;
		18: z3 <= -16'd23;
		19: z3 <= -16'd14;
		20: z3 <= -16'd60;
		21: z3 <= -16'd30;
		22: z3 <= -16'd23;
		23: z3 <= -16'd101;
		24: z3 <= 16'd14;
		25: z3 <= -16'd83;
		26: z3 <= -16'd38;
		27: z3 <= 16'd74;
		28: z3 <= -16'd90;
		29: z3 <= -16'd73;
		30: z3 <= 16'd62;
		31: z3 <= 16'd112;
		32: z3 <= -16'd81;
		33: z3 <= -16'd27;
		34: z3 <= 16'd115;
		35: z3 <= 16'd116;
		36: z3 <= 16'd76;
		37: z3 <= -16'd127;
		38: z3 <= -16'd96;
		39: z3 <= 16'd81;
		40: z3 <= 16'd108;
		41: z3 <= 16'd5;
		42: z3 <= 16'd71;
		43: z3 <= 16'd68;
		44: z3 <= -16'd32;
		45: z3 <= -16'd34;
		46: z3 <= 16'd4;
		47: z3 <= -16'd6;
		48: z3 <= -16'd87;
		49: z3 <= 16'd109;
		50: z3 <= 16'd108;
		51: z3 <= -16'd19;
		52: z3 <= -16'd49;
		53: z3 <= -16'd42;
		54: z3 <= 16'd8;
		55: z3 <= 16'd93;
		56: z3 <= 16'd3;
		57: z3 <= 16'd98;
		58: z3 <= 16'd40;
		59: z3 <= 16'd41;
		60: z3 <= -16'd103;
		61: z3 <= -16'd26;
		62: z3 <= 16'd25;
		63: z3 <= -16'd56;
		64: z3 <= 16'd75;
		65: z3 <= 16'd12;
		66: z3 <= -16'd68;
		67: z3 <= 16'd23;
		68: z3 <= 16'd13;
		69: z3 <= -16'd36;
		70: z3 <= -16'd24;
		71: z3 <= -16'd6;
		72: z3 <= 16'd98;
		73: z3 <= -16'd81;
		74: z3 <= -16'd66;
		75: z3 <= -16'd62;
		76: z3 <= 16'd14;
		77: z3 <= 16'd67;
		78: z3 <= 16'd60;
		79: z3 <= 16'd55;
		80: z3 <= 16'd48;
		81: z3 <= 16'd41;
		82: z3 <= -16'd92;
		83: z3 <= -16'd128;
		84: z3 <= 16'd127;
		85: z3 <= 16'd45;
		86: z3 <= 16'd93;
		87: z3 <= 16'd2;
		88: z3 <= 16'd15;
		89: z3 <= 16'd5;
		90: z3 <= -16'd85;
		91: z3 <= 16'd41;
		92: z3 <= 16'd107;
		93: z3 <= 16'd68;
		94: z3 <= 16'd113;
		95: z3 <= 16'd55;
		96: z3 <= -16'd48;
		97: z3 <= -16'd82;
		98: z3 <= -16'd50;
		99: z3 <= 16'd94;
		100: z3 <= 16'd10;
		101: z3 <= 16'd55;
		102: z3 <= -16'd40;
		103: z3 <= -16'd20;
		104: z3 <= 16'd102;
		105: z3 <= 16'd22;
		106: z3 <= 16'd47;
		107: z3 <= -16'd12;
		108: z3 <= -16'd39;
		109: z3 <= -16'd21;
		110: z3 <= -16'd85;
		111: z3 <= -16'd118;
		112: z3 <= -16'd108;
		113: z3 <= -16'd48;
		114: z3 <= -16'd118;
		115: z3 <= -16'd109;
		116: z3 <= 16'd125;
		117: z3 <= 16'd103;
		118: z3 <= 16'd21;
		119: z3 <= 16'd12;
		120: z3 <= -16'd19;
		121: z3 <= 16'd64;
		122: z3 <= -16'd75;
		123: z3 <= -16'd40;
		124: z3 <= 16'd4;
		125: z3 <= -16'd89;
		126: z3 <= -16'd113;
		127: z3 <= 16'd85;
		endcase
		case(addr4)
		0: z4 <= 16'd74;
		1: z4 <= 16'd120;
		2: z4 <= 16'd39;
		3: z4 <= -16'd125;
		4: z4 <= 16'd69;
		5: z4 <= -16'd26;
		6: z4 <= -16'd115;
		7: z4 <= -16'd84;
		8: z4 <= -16'd123;
		9: z4 <= 16'd107;
		10: z4 <= -16'd27;
		11: z4 <= 16'd118;
		12: z4 <= 16'd88;
		13: z4 <= 16'd91;
		14: z4 <= 16'd23;
		15: z4 <= 16'd64;
		16: z4 <= -16'd103;
		17: z4 <= 16'd74;
		18: z4 <= -16'd23;
		19: z4 <= -16'd14;
		20: z4 <= -16'd60;
		21: z4 <= -16'd30;
		22: z4 <= -16'd23;
		23: z4 <= -16'd101;
		24: z4 <= 16'd14;
		25: z4 <= -16'd83;
		26: z4 <= -16'd38;
		27: z4 <= 16'd74;
		28: z4 <= -16'd90;
		29: z4 <= -16'd73;
		30: z4 <= 16'd62;
		31: z4 <= 16'd112;
		32: z4 <= -16'd81;
		33: z4 <= -16'd27;
		34: z4 <= 16'd115;
		35: z4 <= 16'd116;
		36: z4 <= 16'd76;
		37: z4 <= -16'd127;
		38: z4 <= -16'd96;
		39: z4 <= 16'd81;
		40: z4 <= 16'd108;
		41: z4 <= 16'd5;
		42: z4 <= 16'd71;
		43: z4 <= 16'd68;
		44: z4 <= -16'd32;
		45: z4 <= -16'd34;
		46: z4 <= 16'd4;
		47: z4 <= -16'd6;
		48: z4 <= -16'd87;
		49: z4 <= 16'd109;
		50: z4 <= 16'd108;
		51: z4 <= -16'd19;
		52: z4 <= -16'd49;
		53: z4 <= -16'd42;
		54: z4 <= 16'd8;
		55: z4 <= 16'd93;
		56: z4 <= 16'd3;
		57: z4 <= 16'd98;
		58: z4 <= 16'd40;
		59: z4 <= 16'd41;
		60: z4 <= -16'd103;
		61: z4 <= -16'd26;
		62: z4 <= 16'd25;
		63: z4 <= -16'd56;
		64: z4 <= 16'd75;
		65: z4 <= 16'd12;
		66: z4 <= -16'd68;
		67: z4 <= 16'd23;
		68: z4 <= 16'd13;
		69: z4 <= -16'd36;
		70: z4 <= -16'd24;
		71: z4 <= -16'd6;
		72: z4 <= 16'd98;
		73: z4 <= -16'd81;
		74: z4 <= -16'd66;
		75: z4 <= -16'd62;
		76: z4 <= 16'd14;
		77: z4 <= 16'd67;
		78: z4 <= 16'd60;
		79: z4 <= 16'd55;
		80: z4 <= 16'd48;
		81: z4 <= 16'd41;
		82: z4 <= -16'd92;
		83: z4 <= -16'd128;
		84: z4 <= 16'd127;
		85: z4 <= 16'd45;
		86: z4 <= 16'd93;
		87: z4 <= 16'd2;
		88: z4 <= 16'd15;
		89: z4 <= 16'd5;
		90: z4 <= -16'd85;
		91: z4 <= 16'd41;
		92: z4 <= 16'd107;
		93: z4 <= 16'd68;
		94: z4 <= 16'd113;
		95: z4 <= 16'd55;
		96: z4 <= -16'd48;
		97: z4 <= -16'd82;
		98: z4 <= -16'd50;
		99: z4 <= 16'd94;
		100: z4 <= 16'd10;
		101: z4 <= 16'd55;
		102: z4 <= -16'd40;
		103: z4 <= -16'd20;
		104: z4 <= 16'd102;
		105: z4 <= 16'd22;
		106: z4 <= 16'd47;
		107: z4 <= -16'd12;
		108: z4 <= -16'd39;
		109: z4 <= -16'd21;
		110: z4 <= -16'd85;
		111: z4 <= -16'd118;
		112: z4 <= -16'd108;
		113: z4 <= -16'd48;
		114: z4 <= -16'd118;
		115: z4 <= -16'd109;
		116: z4 <= 16'd125;
		117: z4 <= 16'd103;
		118: z4 <= 16'd21;
		119: z4 <= 16'd12;
		120: z4 <= -16'd19;
		121: z4 <= 16'd64;
		122: z4 <= -16'd75;
		123: z4 <= -16'd40;
		124: z4 <= 16'd4;
		125: z4 <= -16'd89;
		126: z4 <= -16'd113;
		127: z4 <= 16'd85;
		endcase
		case(addr5)
		0: z5 <= 16'd74;
		1: z5 <= 16'd120;
		2: z5 <= 16'd39;
		3: z5 <= -16'd125;
		4: z5 <= 16'd69;
		5: z5 <= -16'd26;
		6: z5 <= -16'd115;
		7: z5 <= -16'd84;
		8: z5 <= -16'd123;
		9: z5 <= 16'd107;
		10: z5 <= -16'd27;
		11: z5 <= 16'd118;
		12: z5 <= 16'd88;
		13: z5 <= 16'd91;
		14: z5 <= 16'd23;
		15: z5 <= 16'd64;
		16: z5 <= -16'd103;
		17: z5 <= 16'd74;
		18: z5 <= -16'd23;
		19: z5 <= -16'd14;
		20: z5 <= -16'd60;
		21: z5 <= -16'd30;
		22: z5 <= -16'd23;
		23: z5 <= -16'd101;
		24: z5 <= 16'd14;
		25: z5 <= -16'd83;
		26: z5 <= -16'd38;
		27: z5 <= 16'd74;
		28: z5 <= -16'd90;
		29: z5 <= -16'd73;
		30: z5 <= 16'd62;
		31: z5 <= 16'd112;
		32: z5 <= -16'd81;
		33: z5 <= -16'd27;
		34: z5 <= 16'd115;
		35: z5 <= 16'd116;
		36: z5 <= 16'd76;
		37: z5 <= -16'd127;
		38: z5 <= -16'd96;
		39: z5 <= 16'd81;
		40: z5 <= 16'd108;
		41: z5 <= 16'd5;
		42: z5 <= 16'd71;
		43: z5 <= 16'd68;
		44: z5 <= -16'd32;
		45: z5 <= -16'd34;
		46: z5 <= 16'd4;
		47: z5 <= -16'd6;
		48: z5 <= -16'd87;
		49: z5 <= 16'd109;
		50: z5 <= 16'd108;
		51: z5 <= -16'd19;
		52: z5 <= -16'd49;
		53: z5 <= -16'd42;
		54: z5 <= 16'd8;
		55: z5 <= 16'd93;
		56: z5 <= 16'd3;
		57: z5 <= 16'd98;
		58: z5 <= 16'd40;
		59: z5 <= 16'd41;
		60: z5 <= -16'd103;
		61: z5 <= -16'd26;
		62: z5 <= 16'd25;
		63: z5 <= -16'd56;
		64: z5 <= 16'd75;
		65: z5 <= 16'd12;
		66: z5 <= -16'd68;
		67: z5 <= 16'd23;
		68: z5 <= 16'd13;
		69: z5 <= -16'd36;
		70: z5 <= -16'd24;
		71: z5 <= -16'd6;
		72: z5 <= 16'd98;
		73: z5 <= -16'd81;
		74: z5 <= -16'd66;
		75: z5 <= -16'd62;
		76: z5 <= 16'd14;
		77: z5 <= 16'd67;
		78: z5 <= 16'd60;
		79: z5 <= 16'd55;
		80: z5 <= 16'd48;
		81: z5 <= 16'd41;
		82: z5 <= -16'd92;
		83: z5 <= -16'd128;
		84: z5 <= 16'd127;
		85: z5 <= 16'd45;
		86: z5 <= 16'd93;
		87: z5 <= 16'd2;
		88: z5 <= 16'd15;
		89: z5 <= 16'd5;
		90: z5 <= -16'd85;
		91: z5 <= 16'd41;
		92: z5 <= 16'd107;
		93: z5 <= 16'd68;
		94: z5 <= 16'd113;
		95: z5 <= 16'd55;
		96: z5 <= -16'd48;
		97: z5 <= -16'd82;
		98: z5 <= -16'd50;
		99: z5 <= 16'd94;
		100: z5 <= 16'd10;
		101: z5 <= 16'd55;
		102: z5 <= -16'd40;
		103: z5 <= -16'd20;
		104: z5 <= 16'd102;
		105: z5 <= 16'd22;
		106: z5 <= 16'd47;
		107: z5 <= -16'd12;
		108: z5 <= -16'd39;
		109: z5 <= -16'd21;
		110: z5 <= -16'd85;
		111: z5 <= -16'd118;
		112: z5 <= -16'd108;
		113: z5 <= -16'd48;
		114: z5 <= -16'd118;
		115: z5 <= -16'd109;
		116: z5 <= 16'd125;
		117: z5 <= 16'd103;
		118: z5 <= 16'd21;
		119: z5 <= 16'd12;
		120: z5 <= -16'd19;
		121: z5 <= 16'd64;
		122: z5 <= -16'd75;
		123: z5 <= -16'd40;
		124: z5 <= 16'd4;
		125: z5 <= -16'd89;
		126: z5 <= -16'd113;
		127: z5 <= 16'd85;
		endcase
		case(addr6)
		0: z6 <= 16'd74;
		1: z6 <= 16'd120;
		2: z6 <= 16'd39;
		3: z6 <= -16'd125;
		4: z6 <= 16'd69;
		5: z6 <= -16'd26;
		6: z6 <= -16'd115;
		7: z6 <= -16'd84;
		8: z6 <= -16'd123;
		9: z6 <= 16'd107;
		10: z6 <= -16'd27;
		11: z6 <= 16'd118;
		12: z6 <= 16'd88;
		13: z6 <= 16'd91;
		14: z6 <= 16'd23;
		15: z6 <= 16'd64;
		16: z6 <= -16'd103;
		17: z6 <= 16'd74;
		18: z6 <= -16'd23;
		19: z6 <= -16'd14;
		20: z6 <= -16'd60;
		21: z6 <= -16'd30;
		22: z6 <= -16'd23;
		23: z6 <= -16'd101;
		24: z6 <= 16'd14;
		25: z6 <= -16'd83;
		26: z6 <= -16'd38;
		27: z6 <= 16'd74;
		28: z6 <= -16'd90;
		29: z6 <= -16'd73;
		30: z6 <= 16'd62;
		31: z6 <= 16'd112;
		32: z6 <= -16'd81;
		33: z6 <= -16'd27;
		34: z6 <= 16'd115;
		35: z6 <= 16'd116;
		36: z6 <= 16'd76;
		37: z6 <= -16'd127;
		38: z6 <= -16'd96;
		39: z6 <= 16'd81;
		40: z6 <= 16'd108;
		41: z6 <= 16'd5;
		42: z6 <= 16'd71;
		43: z6 <= 16'd68;
		44: z6 <= -16'd32;
		45: z6 <= -16'd34;
		46: z6 <= 16'd4;
		47: z6 <= -16'd6;
		48: z6 <= -16'd87;
		49: z6 <= 16'd109;
		50: z6 <= 16'd108;
		51: z6 <= -16'd19;
		52: z6 <= -16'd49;
		53: z6 <= -16'd42;
		54: z6 <= 16'd8;
		55: z6 <= 16'd93;
		56: z6 <= 16'd3;
		57: z6 <= 16'd98;
		58: z6 <= 16'd40;
		59: z6 <= 16'd41;
		60: z6 <= -16'd103;
		61: z6 <= -16'd26;
		62: z6 <= 16'd25;
		63: z6 <= -16'd56;
		64: z6 <= 16'd75;
		65: z6 <= 16'd12;
		66: z6 <= -16'd68;
		67: z6 <= 16'd23;
		68: z6 <= 16'd13;
		69: z6 <= -16'd36;
		70: z6 <= -16'd24;
		71: z6 <= -16'd6;
		72: z6 <= 16'd98;
		73: z6 <= -16'd81;
		74: z6 <= -16'd66;
		75: z6 <= -16'd62;
		76: z6 <= 16'd14;
		77: z6 <= 16'd67;
		78: z6 <= 16'd60;
		79: z6 <= 16'd55;
		80: z6 <= 16'd48;
		81: z6 <= 16'd41;
		82: z6 <= -16'd92;
		83: z6 <= -16'd128;
		84: z6 <= 16'd127;
		85: z6 <= 16'd45;
		86: z6 <= 16'd93;
		87: z6 <= 16'd2;
		88: z6 <= 16'd15;
		89: z6 <= 16'd5;
		90: z6 <= -16'd85;
		91: z6 <= 16'd41;
		92: z6 <= 16'd107;
		93: z6 <= 16'd68;
		94: z6 <= 16'd113;
		95: z6 <= 16'd55;
		96: z6 <= -16'd48;
		97: z6 <= -16'd82;
		98: z6 <= -16'd50;
		99: z6 <= 16'd94;
		100: z6 <= 16'd10;
		101: z6 <= 16'd55;
		102: z6 <= -16'd40;
		103: z6 <= -16'd20;
		104: z6 <= 16'd102;
		105: z6 <= 16'd22;
		106: z6 <= 16'd47;
		107: z6 <= -16'd12;
		108: z6 <= -16'd39;
		109: z6 <= -16'd21;
		110: z6 <= -16'd85;
		111: z6 <= -16'd118;
		112: z6 <= -16'd108;
		113: z6 <= -16'd48;
		114: z6 <= -16'd118;
		115: z6 <= -16'd109;
		116: z6 <= 16'd125;
		117: z6 <= 16'd103;
		118: z6 <= 16'd21;
		119: z6 <= 16'd12;
		120: z6 <= -16'd19;
		121: z6 <= 16'd64;
		122: z6 <= -16'd75;
		123: z6 <= -16'd40;
		124: z6 <= 16'd4;
		125: z6 <= -16'd89;
		126: z6 <= -16'd113;
		127: z6 <= 16'd85;
		endcase
		case(addr7)
		0: z7 <= 16'd74;
		1: z7 <= 16'd120;
		2: z7 <= 16'd39;
		3: z7 <= -16'd125;
		4: z7 <= 16'd69;
		5: z7 <= -16'd26;
		6: z7 <= -16'd115;
		7: z7 <= -16'd84;
		8: z7 <= -16'd123;
		9: z7 <= 16'd107;
		10: z7 <= -16'd27;
		11: z7 <= 16'd118;
		12: z7 <= 16'd88;
		13: z7 <= 16'd91;
		14: z7 <= 16'd23;
		15: z7 <= 16'd64;
		16: z7 <= -16'd103;
		17: z7 <= 16'd74;
		18: z7 <= -16'd23;
		19: z7 <= -16'd14;
		20: z7 <= -16'd60;
		21: z7 <= -16'd30;
		22: z7 <= -16'd23;
		23: z7 <= -16'd101;
		24: z7 <= 16'd14;
		25: z7 <= -16'd83;
		26: z7 <= -16'd38;
		27: z7 <= 16'd74;
		28: z7 <= -16'd90;
		29: z7 <= -16'd73;
		30: z7 <= 16'd62;
		31: z7 <= 16'd112;
		32: z7 <= -16'd81;
		33: z7 <= -16'd27;
		34: z7 <= 16'd115;
		35: z7 <= 16'd116;
		36: z7 <= 16'd76;
		37: z7 <= -16'd127;
		38: z7 <= -16'd96;
		39: z7 <= 16'd81;
		40: z7 <= 16'd108;
		41: z7 <= 16'd5;
		42: z7 <= 16'd71;
		43: z7 <= 16'd68;
		44: z7 <= -16'd32;
		45: z7 <= -16'd34;
		46: z7 <= 16'd4;
		47: z7 <= -16'd6;
		48: z7 <= -16'd87;
		49: z7 <= 16'd109;
		50: z7 <= 16'd108;
		51: z7 <= -16'd19;
		52: z7 <= -16'd49;
		53: z7 <= -16'd42;
		54: z7 <= 16'd8;
		55: z7 <= 16'd93;
		56: z7 <= 16'd3;
		57: z7 <= 16'd98;
		58: z7 <= 16'd40;
		59: z7 <= 16'd41;
		60: z7 <= -16'd103;
		61: z7 <= -16'd26;
		62: z7 <= 16'd25;
		63: z7 <= -16'd56;
		64: z7 <= 16'd75;
		65: z7 <= 16'd12;
		66: z7 <= -16'd68;
		67: z7 <= 16'd23;
		68: z7 <= 16'd13;
		69: z7 <= -16'd36;
		70: z7 <= -16'd24;
		71: z7 <= -16'd6;
		72: z7 <= 16'd98;
		73: z7 <= -16'd81;
		74: z7 <= -16'd66;
		75: z7 <= -16'd62;
		76: z7 <= 16'd14;
		77: z7 <= 16'd67;
		78: z7 <= 16'd60;
		79: z7 <= 16'd55;
		80: z7 <= 16'd48;
		81: z7 <= 16'd41;
		82: z7 <= -16'd92;
		83: z7 <= -16'd128;
		84: z7 <= 16'd127;
		85: z7 <= 16'd45;
		86: z7 <= 16'd93;
		87: z7 <= 16'd2;
		88: z7 <= 16'd15;
		89: z7 <= 16'd5;
		90: z7 <= -16'd85;
		91: z7 <= 16'd41;
		92: z7 <= 16'd107;
		93: z7 <= 16'd68;
		94: z7 <= 16'd113;
		95: z7 <= 16'd55;
		96: z7 <= -16'd48;
		97: z7 <= -16'd82;
		98: z7 <= -16'd50;
		99: z7 <= 16'd94;
		100: z7 <= 16'd10;
		101: z7 <= 16'd55;
		102: z7 <= -16'd40;
		103: z7 <= -16'd20;
		104: z7 <= 16'd102;
		105: z7 <= 16'd22;
		106: z7 <= 16'd47;
		107: z7 <= -16'd12;
		108: z7 <= -16'd39;
		109: z7 <= -16'd21;
		110: z7 <= -16'd85;
		111: z7 <= -16'd118;
		112: z7 <= -16'd108;
		113: z7 <= -16'd48;
		114: z7 <= -16'd118;
		115: z7 <= -16'd109;
		116: z7 <= 16'd125;
		117: z7 <= 16'd103;
		118: z7 <= 16'd21;
		119: z7 <= 16'd12;
		120: z7 <= -16'd19;
		121: z7 <= 16'd64;
		122: z7 <= -16'd75;
		123: z7 <= -16'd40;
		124: z7 <= 16'd4;
		125: z7 <= -16'd89;
		126: z7 <= -16'd113;
		127: z7 <= 16'd85;
		endcase
		case(addr8)
		0: z8 <= 16'd74;
		1: z8 <= 16'd120;
		2: z8 <= 16'd39;
		3: z8 <= -16'd125;
		4: z8 <= 16'd69;
		5: z8 <= -16'd26;
		6: z8 <= -16'd115;
		7: z8 <= -16'd84;
		8: z8 <= -16'd123;
		9: z8 <= 16'd107;
		10: z8 <= -16'd27;
		11: z8 <= 16'd118;
		12: z8 <= 16'd88;
		13: z8 <= 16'd91;
		14: z8 <= 16'd23;
		15: z8 <= 16'd64;
		16: z8 <= -16'd103;
		17: z8 <= 16'd74;
		18: z8 <= -16'd23;
		19: z8 <= -16'd14;
		20: z8 <= -16'd60;
		21: z8 <= -16'd30;
		22: z8 <= -16'd23;
		23: z8 <= -16'd101;
		24: z8 <= 16'd14;
		25: z8 <= -16'd83;
		26: z8 <= -16'd38;
		27: z8 <= 16'd74;
		28: z8 <= -16'd90;
		29: z8 <= -16'd73;
		30: z8 <= 16'd62;
		31: z8 <= 16'd112;
		32: z8 <= -16'd81;
		33: z8 <= -16'd27;
		34: z8 <= 16'd115;
		35: z8 <= 16'd116;
		36: z8 <= 16'd76;
		37: z8 <= -16'd127;
		38: z8 <= -16'd96;
		39: z8 <= 16'd81;
		40: z8 <= 16'd108;
		41: z8 <= 16'd5;
		42: z8 <= 16'd71;
		43: z8 <= 16'd68;
		44: z8 <= -16'd32;
		45: z8 <= -16'd34;
		46: z8 <= 16'd4;
		47: z8 <= -16'd6;
		48: z8 <= -16'd87;
		49: z8 <= 16'd109;
		50: z8 <= 16'd108;
		51: z8 <= -16'd19;
		52: z8 <= -16'd49;
		53: z8 <= -16'd42;
		54: z8 <= 16'd8;
		55: z8 <= 16'd93;
		56: z8 <= 16'd3;
		57: z8 <= 16'd98;
		58: z8 <= 16'd40;
		59: z8 <= 16'd41;
		60: z8 <= -16'd103;
		61: z8 <= -16'd26;
		62: z8 <= 16'd25;
		63: z8 <= -16'd56;
		64: z8 <= 16'd75;
		65: z8 <= 16'd12;
		66: z8 <= -16'd68;
		67: z8 <= 16'd23;
		68: z8 <= 16'd13;
		69: z8 <= -16'd36;
		70: z8 <= -16'd24;
		71: z8 <= -16'd6;
		72: z8 <= 16'd98;
		73: z8 <= -16'd81;
		74: z8 <= -16'd66;
		75: z8 <= -16'd62;
		76: z8 <= 16'd14;
		77: z8 <= 16'd67;
		78: z8 <= 16'd60;
		79: z8 <= 16'd55;
		80: z8 <= 16'd48;
		81: z8 <= 16'd41;
		82: z8 <= -16'd92;
		83: z8 <= -16'd128;
		84: z8 <= 16'd127;
		85: z8 <= 16'd45;
		86: z8 <= 16'd93;
		87: z8 <= 16'd2;
		88: z8 <= 16'd15;
		89: z8 <= 16'd5;
		90: z8 <= -16'd85;
		91: z8 <= 16'd41;
		92: z8 <= 16'd107;
		93: z8 <= 16'd68;
		94: z8 <= 16'd113;
		95: z8 <= 16'd55;
		96: z8 <= -16'd48;
		97: z8 <= -16'd82;
		98: z8 <= -16'd50;
		99: z8 <= 16'd94;
		100: z8 <= 16'd10;
		101: z8 <= 16'd55;
		102: z8 <= -16'd40;
		103: z8 <= -16'd20;
		104: z8 <= 16'd102;
		105: z8 <= 16'd22;
		106: z8 <= 16'd47;
		107: z8 <= -16'd12;
		108: z8 <= -16'd39;
		109: z8 <= -16'd21;
		110: z8 <= -16'd85;
		111: z8 <= -16'd118;
		112: z8 <= -16'd108;
		113: z8 <= -16'd48;
		114: z8 <= -16'd118;
		115: z8 <= -16'd109;
		116: z8 <= 16'd125;
		117: z8 <= 16'd103;
		118: z8 <= 16'd21;
		119: z8 <= 16'd12;
		120: z8 <= -16'd19;
		121: z8 <= 16'd64;
		122: z8 <= -16'd75;
		123: z8 <= -16'd40;
		124: z8 <= 16'd4;
		125: z8 <= -16'd89;
		126: z8 <= -16'd113;
		127: z8 <= 16'd85;
		endcase
		case(addr9)
		0: z9 <= 16'd74;
		1: z9 <= 16'd120;
		2: z9 <= 16'd39;
		3: z9 <= -16'd125;
		4: z9 <= 16'd69;
		5: z9 <= -16'd26;
		6: z9 <= -16'd115;
		7: z9 <= -16'd84;
		8: z9 <= -16'd123;
		9: z9 <= 16'd107;
		10: z9 <= -16'd27;
		11: z9 <= 16'd118;
		12: z9 <= 16'd88;
		13: z9 <= 16'd91;
		14: z9 <= 16'd23;
		15: z9 <= 16'd64;
		16: z9 <= -16'd103;
		17: z9 <= 16'd74;
		18: z9 <= -16'd23;
		19: z9 <= -16'd14;
		20: z9 <= -16'd60;
		21: z9 <= -16'd30;
		22: z9 <= -16'd23;
		23: z9 <= -16'd101;
		24: z9 <= 16'd14;
		25: z9 <= -16'd83;
		26: z9 <= -16'd38;
		27: z9 <= 16'd74;
		28: z9 <= -16'd90;
		29: z9 <= -16'd73;
		30: z9 <= 16'd62;
		31: z9 <= 16'd112;
		32: z9 <= -16'd81;
		33: z9 <= -16'd27;
		34: z9 <= 16'd115;
		35: z9 <= 16'd116;
		36: z9 <= 16'd76;
		37: z9 <= -16'd127;
		38: z9 <= -16'd96;
		39: z9 <= 16'd81;
		40: z9 <= 16'd108;
		41: z9 <= 16'd5;
		42: z9 <= 16'd71;
		43: z9 <= 16'd68;
		44: z9 <= -16'd32;
		45: z9 <= -16'd34;
		46: z9 <= 16'd4;
		47: z9 <= -16'd6;
		48: z9 <= -16'd87;
		49: z9 <= 16'd109;
		50: z9 <= 16'd108;
		51: z9 <= -16'd19;
		52: z9 <= -16'd49;
		53: z9 <= -16'd42;
		54: z9 <= 16'd8;
		55: z9 <= 16'd93;
		56: z9 <= 16'd3;
		57: z9 <= 16'd98;
		58: z9 <= 16'd40;
		59: z9 <= 16'd41;
		60: z9 <= -16'd103;
		61: z9 <= -16'd26;
		62: z9 <= 16'd25;
		63: z9 <= -16'd56;
		64: z9 <= 16'd75;
		65: z9 <= 16'd12;
		66: z9 <= -16'd68;
		67: z9 <= 16'd23;
		68: z9 <= 16'd13;
		69: z9 <= -16'd36;
		70: z9 <= -16'd24;
		71: z9 <= -16'd6;
		72: z9 <= 16'd98;
		73: z9 <= -16'd81;
		74: z9 <= -16'd66;
		75: z9 <= -16'd62;
		76: z9 <= 16'd14;
		77: z9 <= 16'd67;
		78: z9 <= 16'd60;
		79: z9 <= 16'd55;
		80: z9 <= 16'd48;
		81: z9 <= 16'd41;
		82: z9 <= -16'd92;
		83: z9 <= -16'd128;
		84: z9 <= 16'd127;
		85: z9 <= 16'd45;
		86: z9 <= 16'd93;
		87: z9 <= 16'd2;
		88: z9 <= 16'd15;
		89: z9 <= 16'd5;
		90: z9 <= -16'd85;
		91: z9 <= 16'd41;
		92: z9 <= 16'd107;
		93: z9 <= 16'd68;
		94: z9 <= 16'd113;
		95: z9 <= 16'd55;
		96: z9 <= -16'd48;
		97: z9 <= -16'd82;
		98: z9 <= -16'd50;
		99: z9 <= 16'd94;
		100: z9 <= 16'd10;
		101: z9 <= 16'd55;
		102: z9 <= -16'd40;
		103: z9 <= -16'd20;
		104: z9 <= 16'd102;
		105: z9 <= 16'd22;
		106: z9 <= 16'd47;
		107: z9 <= -16'd12;
		108: z9 <= -16'd39;
		109: z9 <= -16'd21;
		110: z9 <= -16'd85;
		111: z9 <= -16'd118;
		112: z9 <= -16'd108;
		113: z9 <= -16'd48;
		114: z9 <= -16'd118;
		115: z9 <= -16'd109;
		116: z9 <= 16'd125;
		117: z9 <= 16'd103;
		118: z9 <= 16'd21;
		119: z9 <= 16'd12;
		120: z9 <= -16'd19;
		121: z9 <= 16'd64;
		122: z9 <= -16'd75;
		123: z9 <= -16'd40;
		124: z9 <= 16'd4;
		125: z9 <= -16'd89;
		126: z9 <= -16'd113;
		127: z9 <= 16'd85;
		endcase
		case(addr10)
		0: z10 <= 16'd74;
		1: z10 <= 16'd120;
		2: z10 <= 16'd39;
		3: z10 <= -16'd125;
		4: z10 <= 16'd69;
		5: z10 <= -16'd26;
		6: z10 <= -16'd115;
		7: z10 <= -16'd84;
		8: z10 <= -16'd123;
		9: z10 <= 16'd107;
		10: z10 <= -16'd27;
		11: z10 <= 16'd118;
		12: z10 <= 16'd88;
		13: z10 <= 16'd91;
		14: z10 <= 16'd23;
		15: z10 <= 16'd64;
		16: z10 <= -16'd103;
		17: z10 <= 16'd74;
		18: z10 <= -16'd23;
		19: z10 <= -16'd14;
		20: z10 <= -16'd60;
		21: z10 <= -16'd30;
		22: z10 <= -16'd23;
		23: z10 <= -16'd101;
		24: z10 <= 16'd14;
		25: z10 <= -16'd83;
		26: z10 <= -16'd38;
		27: z10 <= 16'd74;
		28: z10 <= -16'd90;
		29: z10 <= -16'd73;
		30: z10 <= 16'd62;
		31: z10 <= 16'd112;
		32: z10 <= -16'd81;
		33: z10 <= -16'd27;
		34: z10 <= 16'd115;
		35: z10 <= 16'd116;
		36: z10 <= 16'd76;
		37: z10 <= -16'd127;
		38: z10 <= -16'd96;
		39: z10 <= 16'd81;
		40: z10 <= 16'd108;
		41: z10 <= 16'd5;
		42: z10 <= 16'd71;
		43: z10 <= 16'd68;
		44: z10 <= -16'd32;
		45: z10 <= -16'd34;
		46: z10 <= 16'd4;
		47: z10 <= -16'd6;
		48: z10 <= -16'd87;
		49: z10 <= 16'd109;
		50: z10 <= 16'd108;
		51: z10 <= -16'd19;
		52: z10 <= -16'd49;
		53: z10 <= -16'd42;
		54: z10 <= 16'd8;
		55: z10 <= 16'd93;
		56: z10 <= 16'd3;
		57: z10 <= 16'd98;
		58: z10 <= 16'd40;
		59: z10 <= 16'd41;
		60: z10 <= -16'd103;
		61: z10 <= -16'd26;
		62: z10 <= 16'd25;
		63: z10 <= -16'd56;
		64: z10 <= 16'd75;
		65: z10 <= 16'd12;
		66: z10 <= -16'd68;
		67: z10 <= 16'd23;
		68: z10 <= 16'd13;
		69: z10 <= -16'd36;
		70: z10 <= -16'd24;
		71: z10 <= -16'd6;
		72: z10 <= 16'd98;
		73: z10 <= -16'd81;
		74: z10 <= -16'd66;
		75: z10 <= -16'd62;
		76: z10 <= 16'd14;
		77: z10 <= 16'd67;
		78: z10 <= 16'd60;
		79: z10 <= 16'd55;
		80: z10 <= 16'd48;
		81: z10 <= 16'd41;
		82: z10 <= -16'd92;
		83: z10 <= -16'd128;
		84: z10 <= 16'd127;
		85: z10 <= 16'd45;
		86: z10 <= 16'd93;
		87: z10 <= 16'd2;
		88: z10 <= 16'd15;
		89: z10 <= 16'd5;
		90: z10 <= -16'd85;
		91: z10 <= 16'd41;
		92: z10 <= 16'd107;
		93: z10 <= 16'd68;
		94: z10 <= 16'd113;
		95: z10 <= 16'd55;
		96: z10 <= -16'd48;
		97: z10 <= -16'd82;
		98: z10 <= -16'd50;
		99: z10 <= 16'd94;
		100: z10 <= 16'd10;
		101: z10 <= 16'd55;
		102: z10 <= -16'd40;
		103: z10 <= -16'd20;
		104: z10 <= 16'd102;
		105: z10 <= 16'd22;
		106: z10 <= 16'd47;
		107: z10 <= -16'd12;
		108: z10 <= -16'd39;
		109: z10 <= -16'd21;
		110: z10 <= -16'd85;
		111: z10 <= -16'd118;
		112: z10 <= -16'd108;
		113: z10 <= -16'd48;
		114: z10 <= -16'd118;
		115: z10 <= -16'd109;
		116: z10 <= 16'd125;
		117: z10 <= 16'd103;
		118: z10 <= 16'd21;
		119: z10 <= 16'd12;
		120: z10 <= -16'd19;
		121: z10 <= 16'd64;
		122: z10 <= -16'd75;
		123: z10 <= -16'd40;
		124: z10 <= 16'd4;
		125: z10 <= -16'd89;
		126: z10 <= -16'd113;
		127: z10 <= 16'd85;
		endcase
		case(addr11)
		0: z11 <= 16'd74;
		1: z11 <= 16'd120;
		2: z11 <= 16'd39;
		3: z11 <= -16'd125;
		4: z11 <= 16'd69;
		5: z11 <= -16'd26;
		6: z11 <= -16'd115;
		7: z11 <= -16'd84;
		8: z11 <= -16'd123;
		9: z11 <= 16'd107;
		10: z11 <= -16'd27;
		11: z11 <= 16'd118;
		12: z11 <= 16'd88;
		13: z11 <= 16'd91;
		14: z11 <= 16'd23;
		15: z11 <= 16'd64;
		16: z11 <= -16'd103;
		17: z11 <= 16'd74;
		18: z11 <= -16'd23;
		19: z11 <= -16'd14;
		20: z11 <= -16'd60;
		21: z11 <= -16'd30;
		22: z11 <= -16'd23;
		23: z11 <= -16'd101;
		24: z11 <= 16'd14;
		25: z11 <= -16'd83;
		26: z11 <= -16'd38;
		27: z11 <= 16'd74;
		28: z11 <= -16'd90;
		29: z11 <= -16'd73;
		30: z11 <= 16'd62;
		31: z11 <= 16'd112;
		32: z11 <= -16'd81;
		33: z11 <= -16'd27;
		34: z11 <= 16'd115;
		35: z11 <= 16'd116;
		36: z11 <= 16'd76;
		37: z11 <= -16'd127;
		38: z11 <= -16'd96;
		39: z11 <= 16'd81;
		40: z11 <= 16'd108;
		41: z11 <= 16'd5;
		42: z11 <= 16'd71;
		43: z11 <= 16'd68;
		44: z11 <= -16'd32;
		45: z11 <= -16'd34;
		46: z11 <= 16'd4;
		47: z11 <= -16'd6;
		48: z11 <= -16'd87;
		49: z11 <= 16'd109;
		50: z11 <= 16'd108;
		51: z11 <= -16'd19;
		52: z11 <= -16'd49;
		53: z11 <= -16'd42;
		54: z11 <= 16'd8;
		55: z11 <= 16'd93;
		56: z11 <= 16'd3;
		57: z11 <= 16'd98;
		58: z11 <= 16'd40;
		59: z11 <= 16'd41;
		60: z11 <= -16'd103;
		61: z11 <= -16'd26;
		62: z11 <= 16'd25;
		63: z11 <= -16'd56;
		64: z11 <= 16'd75;
		65: z11 <= 16'd12;
		66: z11 <= -16'd68;
		67: z11 <= 16'd23;
		68: z11 <= 16'd13;
		69: z11 <= -16'd36;
		70: z11 <= -16'd24;
		71: z11 <= -16'd6;
		72: z11 <= 16'd98;
		73: z11 <= -16'd81;
		74: z11 <= -16'd66;
		75: z11 <= -16'd62;
		76: z11 <= 16'd14;
		77: z11 <= 16'd67;
		78: z11 <= 16'd60;
		79: z11 <= 16'd55;
		80: z11 <= 16'd48;
		81: z11 <= 16'd41;
		82: z11 <= -16'd92;
		83: z11 <= -16'd128;
		84: z11 <= 16'd127;
		85: z11 <= 16'd45;
		86: z11 <= 16'd93;
		87: z11 <= 16'd2;
		88: z11 <= 16'd15;
		89: z11 <= 16'd5;
		90: z11 <= -16'd85;
		91: z11 <= 16'd41;
		92: z11 <= 16'd107;
		93: z11 <= 16'd68;
		94: z11 <= 16'd113;
		95: z11 <= 16'd55;
		96: z11 <= -16'd48;
		97: z11 <= -16'd82;
		98: z11 <= -16'd50;
		99: z11 <= 16'd94;
		100: z11 <= 16'd10;
		101: z11 <= 16'd55;
		102: z11 <= -16'd40;
		103: z11 <= -16'd20;
		104: z11 <= 16'd102;
		105: z11 <= 16'd22;
		106: z11 <= 16'd47;
		107: z11 <= -16'd12;
		108: z11 <= -16'd39;
		109: z11 <= -16'd21;
		110: z11 <= -16'd85;
		111: z11 <= -16'd118;
		112: z11 <= -16'd108;
		113: z11 <= -16'd48;
		114: z11 <= -16'd118;
		115: z11 <= -16'd109;
		116: z11 <= 16'd125;
		117: z11 <= 16'd103;
		118: z11 <= 16'd21;
		119: z11 <= 16'd12;
		120: z11 <= -16'd19;
		121: z11 <= 16'd64;
		122: z11 <= -16'd75;
		123: z11 <= -16'd40;
		124: z11 <= 16'd4;
		125: z11 <= -16'd89;
		126: z11 <= -16'd113;
		127: z11 <= 16'd85;
		endcase
		case(addr12)
		0: z12 <= 16'd74;
		1: z12 <= 16'd120;
		2: z12 <= 16'd39;
		3: z12 <= -16'd125;
		4: z12 <= 16'd69;
		5: z12 <= -16'd26;
		6: z12 <= -16'd115;
		7: z12 <= -16'd84;
		8: z12 <= -16'd123;
		9: z12 <= 16'd107;
		10: z12 <= -16'd27;
		11: z12 <= 16'd118;
		12: z12 <= 16'd88;
		13: z12 <= 16'd91;
		14: z12 <= 16'd23;
		15: z12 <= 16'd64;
		16: z12 <= -16'd103;
		17: z12 <= 16'd74;
		18: z12 <= -16'd23;
		19: z12 <= -16'd14;
		20: z12 <= -16'd60;
		21: z12 <= -16'd30;
		22: z12 <= -16'd23;
		23: z12 <= -16'd101;
		24: z12 <= 16'd14;
		25: z12 <= -16'd83;
		26: z12 <= -16'd38;
		27: z12 <= 16'd74;
		28: z12 <= -16'd90;
		29: z12 <= -16'd73;
		30: z12 <= 16'd62;
		31: z12 <= 16'd112;
		32: z12 <= -16'd81;
		33: z12 <= -16'd27;
		34: z12 <= 16'd115;
		35: z12 <= 16'd116;
		36: z12 <= 16'd76;
		37: z12 <= -16'd127;
		38: z12 <= -16'd96;
		39: z12 <= 16'd81;
		40: z12 <= 16'd108;
		41: z12 <= 16'd5;
		42: z12 <= 16'd71;
		43: z12 <= 16'd68;
		44: z12 <= -16'd32;
		45: z12 <= -16'd34;
		46: z12 <= 16'd4;
		47: z12 <= -16'd6;
		48: z12 <= -16'd87;
		49: z12 <= 16'd109;
		50: z12 <= 16'd108;
		51: z12 <= -16'd19;
		52: z12 <= -16'd49;
		53: z12 <= -16'd42;
		54: z12 <= 16'd8;
		55: z12 <= 16'd93;
		56: z12 <= 16'd3;
		57: z12 <= 16'd98;
		58: z12 <= 16'd40;
		59: z12 <= 16'd41;
		60: z12 <= -16'd103;
		61: z12 <= -16'd26;
		62: z12 <= 16'd25;
		63: z12 <= -16'd56;
		64: z12 <= 16'd75;
		65: z12 <= 16'd12;
		66: z12 <= -16'd68;
		67: z12 <= 16'd23;
		68: z12 <= 16'd13;
		69: z12 <= -16'd36;
		70: z12 <= -16'd24;
		71: z12 <= -16'd6;
		72: z12 <= 16'd98;
		73: z12 <= -16'd81;
		74: z12 <= -16'd66;
		75: z12 <= -16'd62;
		76: z12 <= 16'd14;
		77: z12 <= 16'd67;
		78: z12 <= 16'd60;
		79: z12 <= 16'd55;
		80: z12 <= 16'd48;
		81: z12 <= 16'd41;
		82: z12 <= -16'd92;
		83: z12 <= -16'd128;
		84: z12 <= 16'd127;
		85: z12 <= 16'd45;
		86: z12 <= 16'd93;
		87: z12 <= 16'd2;
		88: z12 <= 16'd15;
		89: z12 <= 16'd5;
		90: z12 <= -16'd85;
		91: z12 <= 16'd41;
		92: z12 <= 16'd107;
		93: z12 <= 16'd68;
		94: z12 <= 16'd113;
		95: z12 <= 16'd55;
		96: z12 <= -16'd48;
		97: z12 <= -16'd82;
		98: z12 <= -16'd50;
		99: z12 <= 16'd94;
		100: z12 <= 16'd10;
		101: z12 <= 16'd55;
		102: z12 <= -16'd40;
		103: z12 <= -16'd20;
		104: z12 <= 16'd102;
		105: z12 <= 16'd22;
		106: z12 <= 16'd47;
		107: z12 <= -16'd12;
		108: z12 <= -16'd39;
		109: z12 <= -16'd21;
		110: z12 <= -16'd85;
		111: z12 <= -16'd118;
		112: z12 <= -16'd108;
		113: z12 <= -16'd48;
		114: z12 <= -16'd118;
		115: z12 <= -16'd109;
		116: z12 <= 16'd125;
		117: z12 <= 16'd103;
		118: z12 <= 16'd21;
		119: z12 <= 16'd12;
		120: z12 <= -16'd19;
		121: z12 <= 16'd64;
		122: z12 <= -16'd75;
		123: z12 <= -16'd40;
		124: z12 <= 16'd4;
		125: z12 <= -16'd89;
		126: z12 <= -16'd113;
		127: z12 <= 16'd85;
		endcase
		case(addr13)
		0: z13 <= 16'd74;
		1: z13 <= 16'd120;
		2: z13 <= 16'd39;
		3: z13 <= -16'd125;
		4: z13 <= 16'd69;
		5: z13 <= -16'd26;
		6: z13 <= -16'd115;
		7: z13 <= -16'd84;
		8: z13 <= -16'd123;
		9: z13 <= 16'd107;
		10: z13 <= -16'd27;
		11: z13 <= 16'd118;
		12: z13 <= 16'd88;
		13: z13 <= 16'd91;
		14: z13 <= 16'd23;
		15: z13 <= 16'd64;
		16: z13 <= -16'd103;
		17: z13 <= 16'd74;
		18: z13 <= -16'd23;
		19: z13 <= -16'd14;
		20: z13 <= -16'd60;
		21: z13 <= -16'd30;
		22: z13 <= -16'd23;
		23: z13 <= -16'd101;
		24: z13 <= 16'd14;
		25: z13 <= -16'd83;
		26: z13 <= -16'd38;
		27: z13 <= 16'd74;
		28: z13 <= -16'd90;
		29: z13 <= -16'd73;
		30: z13 <= 16'd62;
		31: z13 <= 16'd112;
		32: z13 <= -16'd81;
		33: z13 <= -16'd27;
		34: z13 <= 16'd115;
		35: z13 <= 16'd116;
		36: z13 <= 16'd76;
		37: z13 <= -16'd127;
		38: z13 <= -16'd96;
		39: z13 <= 16'd81;
		40: z13 <= 16'd108;
		41: z13 <= 16'd5;
		42: z13 <= 16'd71;
		43: z13 <= 16'd68;
		44: z13 <= -16'd32;
		45: z13 <= -16'd34;
		46: z13 <= 16'd4;
		47: z13 <= -16'd6;
		48: z13 <= -16'd87;
		49: z13 <= 16'd109;
		50: z13 <= 16'd108;
		51: z13 <= -16'd19;
		52: z13 <= -16'd49;
		53: z13 <= -16'd42;
		54: z13 <= 16'd8;
		55: z13 <= 16'd93;
		56: z13 <= 16'd3;
		57: z13 <= 16'd98;
		58: z13 <= 16'd40;
		59: z13 <= 16'd41;
		60: z13 <= -16'd103;
		61: z13 <= -16'd26;
		62: z13 <= 16'd25;
		63: z13 <= -16'd56;
		64: z13 <= 16'd75;
		65: z13 <= 16'd12;
		66: z13 <= -16'd68;
		67: z13 <= 16'd23;
		68: z13 <= 16'd13;
		69: z13 <= -16'd36;
		70: z13 <= -16'd24;
		71: z13 <= -16'd6;
		72: z13 <= 16'd98;
		73: z13 <= -16'd81;
		74: z13 <= -16'd66;
		75: z13 <= -16'd62;
		76: z13 <= 16'd14;
		77: z13 <= 16'd67;
		78: z13 <= 16'd60;
		79: z13 <= 16'd55;
		80: z13 <= 16'd48;
		81: z13 <= 16'd41;
		82: z13 <= -16'd92;
		83: z13 <= -16'd128;
		84: z13 <= 16'd127;
		85: z13 <= 16'd45;
		86: z13 <= 16'd93;
		87: z13 <= 16'd2;
		88: z13 <= 16'd15;
		89: z13 <= 16'd5;
		90: z13 <= -16'd85;
		91: z13 <= 16'd41;
		92: z13 <= 16'd107;
		93: z13 <= 16'd68;
		94: z13 <= 16'd113;
		95: z13 <= 16'd55;
		96: z13 <= -16'd48;
		97: z13 <= -16'd82;
		98: z13 <= -16'd50;
		99: z13 <= 16'd94;
		100: z13 <= 16'd10;
		101: z13 <= 16'd55;
		102: z13 <= -16'd40;
		103: z13 <= -16'd20;
		104: z13 <= 16'd102;
		105: z13 <= 16'd22;
		106: z13 <= 16'd47;
		107: z13 <= -16'd12;
		108: z13 <= -16'd39;
		109: z13 <= -16'd21;
		110: z13 <= -16'd85;
		111: z13 <= -16'd118;
		112: z13 <= -16'd108;
		113: z13 <= -16'd48;
		114: z13 <= -16'd118;
		115: z13 <= -16'd109;
		116: z13 <= 16'd125;
		117: z13 <= 16'd103;
		118: z13 <= 16'd21;
		119: z13 <= 16'd12;
		120: z13 <= -16'd19;
		121: z13 <= 16'd64;
		122: z13 <= -16'd75;
		123: z13 <= -16'd40;
		124: z13 <= 16'd4;
		125: z13 <= -16'd89;
		126: z13 <= -16'd113;
		127: z13 <= 16'd85;
		endcase
		case(addr14)
		0: z14 <= 16'd74;
		1: z14 <= 16'd120;
		2: z14 <= 16'd39;
		3: z14 <= -16'd125;
		4: z14 <= 16'd69;
		5: z14 <= -16'd26;
		6: z14 <= -16'd115;
		7: z14 <= -16'd84;
		8: z14 <= -16'd123;
		9: z14 <= 16'd107;
		10: z14 <= -16'd27;
		11: z14 <= 16'd118;
		12: z14 <= 16'd88;
		13: z14 <= 16'd91;
		14: z14 <= 16'd23;
		15: z14 <= 16'd64;
		16: z14 <= -16'd103;
		17: z14 <= 16'd74;
		18: z14 <= -16'd23;
		19: z14 <= -16'd14;
		20: z14 <= -16'd60;
		21: z14 <= -16'd30;
		22: z14 <= -16'd23;
		23: z14 <= -16'd101;
		24: z14 <= 16'd14;
		25: z14 <= -16'd83;
		26: z14 <= -16'd38;
		27: z14 <= 16'd74;
		28: z14 <= -16'd90;
		29: z14 <= -16'd73;
		30: z14 <= 16'd62;
		31: z14 <= 16'd112;
		32: z14 <= -16'd81;
		33: z14 <= -16'd27;
		34: z14 <= 16'd115;
		35: z14 <= 16'd116;
		36: z14 <= 16'd76;
		37: z14 <= -16'd127;
		38: z14 <= -16'd96;
		39: z14 <= 16'd81;
		40: z14 <= 16'd108;
		41: z14 <= 16'd5;
		42: z14 <= 16'd71;
		43: z14 <= 16'd68;
		44: z14 <= -16'd32;
		45: z14 <= -16'd34;
		46: z14 <= 16'd4;
		47: z14 <= -16'd6;
		48: z14 <= -16'd87;
		49: z14 <= 16'd109;
		50: z14 <= 16'd108;
		51: z14 <= -16'd19;
		52: z14 <= -16'd49;
		53: z14 <= -16'd42;
		54: z14 <= 16'd8;
		55: z14 <= 16'd93;
		56: z14 <= 16'd3;
		57: z14 <= 16'd98;
		58: z14 <= 16'd40;
		59: z14 <= 16'd41;
		60: z14 <= -16'd103;
		61: z14 <= -16'd26;
		62: z14 <= 16'd25;
		63: z14 <= -16'd56;
		64: z14 <= 16'd75;
		65: z14 <= 16'd12;
		66: z14 <= -16'd68;
		67: z14 <= 16'd23;
		68: z14 <= 16'd13;
		69: z14 <= -16'd36;
		70: z14 <= -16'd24;
		71: z14 <= -16'd6;
		72: z14 <= 16'd98;
		73: z14 <= -16'd81;
		74: z14 <= -16'd66;
		75: z14 <= -16'd62;
		76: z14 <= 16'd14;
		77: z14 <= 16'd67;
		78: z14 <= 16'd60;
		79: z14 <= 16'd55;
		80: z14 <= 16'd48;
		81: z14 <= 16'd41;
		82: z14 <= -16'd92;
		83: z14 <= -16'd128;
		84: z14 <= 16'd127;
		85: z14 <= 16'd45;
		86: z14 <= 16'd93;
		87: z14 <= 16'd2;
		88: z14 <= 16'd15;
		89: z14 <= 16'd5;
		90: z14 <= -16'd85;
		91: z14 <= 16'd41;
		92: z14 <= 16'd107;
		93: z14 <= 16'd68;
		94: z14 <= 16'd113;
		95: z14 <= 16'd55;
		96: z14 <= -16'd48;
		97: z14 <= -16'd82;
		98: z14 <= -16'd50;
		99: z14 <= 16'd94;
		100: z14 <= 16'd10;
		101: z14 <= 16'd55;
		102: z14 <= -16'd40;
		103: z14 <= -16'd20;
		104: z14 <= 16'd102;
		105: z14 <= 16'd22;
		106: z14 <= 16'd47;
		107: z14 <= -16'd12;
		108: z14 <= -16'd39;
		109: z14 <= -16'd21;
		110: z14 <= -16'd85;
		111: z14 <= -16'd118;
		112: z14 <= -16'd108;
		113: z14 <= -16'd48;
		114: z14 <= -16'd118;
		115: z14 <= -16'd109;
		116: z14 <= 16'd125;
		117: z14 <= 16'd103;
		118: z14 <= 16'd21;
		119: z14 <= 16'd12;
		120: z14 <= -16'd19;
		121: z14 <= 16'd64;
		122: z14 <= -16'd75;
		123: z14 <= -16'd40;
		124: z14 <= 16'd4;
		125: z14 <= -16'd89;
		126: z14 <= -16'd113;
		127: z14 <= 16'd85;
		endcase
		case(addr15)
		0: z15 <= 16'd74;
		1: z15 <= 16'd120;
		2: z15 <= 16'd39;
		3: z15 <= -16'd125;
		4: z15 <= 16'd69;
		5: z15 <= -16'd26;
		6: z15 <= -16'd115;
		7: z15 <= -16'd84;
		8: z15 <= -16'd123;
		9: z15 <= 16'd107;
		10: z15 <= -16'd27;
		11: z15 <= 16'd118;
		12: z15 <= 16'd88;
		13: z15 <= 16'd91;
		14: z15 <= 16'd23;
		15: z15 <= 16'd64;
		16: z15 <= -16'd103;
		17: z15 <= 16'd74;
		18: z15 <= -16'd23;
		19: z15 <= -16'd14;
		20: z15 <= -16'd60;
		21: z15 <= -16'd30;
		22: z15 <= -16'd23;
		23: z15 <= -16'd101;
		24: z15 <= 16'd14;
		25: z15 <= -16'd83;
		26: z15 <= -16'd38;
		27: z15 <= 16'd74;
		28: z15 <= -16'd90;
		29: z15 <= -16'd73;
		30: z15 <= 16'd62;
		31: z15 <= 16'd112;
		32: z15 <= -16'd81;
		33: z15 <= -16'd27;
		34: z15 <= 16'd115;
		35: z15 <= 16'd116;
		36: z15 <= 16'd76;
		37: z15 <= -16'd127;
		38: z15 <= -16'd96;
		39: z15 <= 16'd81;
		40: z15 <= 16'd108;
		41: z15 <= 16'd5;
		42: z15 <= 16'd71;
		43: z15 <= 16'd68;
		44: z15 <= -16'd32;
		45: z15 <= -16'd34;
		46: z15 <= 16'd4;
		47: z15 <= -16'd6;
		48: z15 <= -16'd87;
		49: z15 <= 16'd109;
		50: z15 <= 16'd108;
		51: z15 <= -16'd19;
		52: z15 <= -16'd49;
		53: z15 <= -16'd42;
		54: z15 <= 16'd8;
		55: z15 <= 16'd93;
		56: z15 <= 16'd3;
		57: z15 <= 16'd98;
		58: z15 <= 16'd40;
		59: z15 <= 16'd41;
		60: z15 <= -16'd103;
		61: z15 <= -16'd26;
		62: z15 <= 16'd25;
		63: z15 <= -16'd56;
		64: z15 <= 16'd75;
		65: z15 <= 16'd12;
		66: z15 <= -16'd68;
		67: z15 <= 16'd23;
		68: z15 <= 16'd13;
		69: z15 <= -16'd36;
		70: z15 <= -16'd24;
		71: z15 <= -16'd6;
		72: z15 <= 16'd98;
		73: z15 <= -16'd81;
		74: z15 <= -16'd66;
		75: z15 <= -16'd62;
		76: z15 <= 16'd14;
		77: z15 <= 16'd67;
		78: z15 <= 16'd60;
		79: z15 <= 16'd55;
		80: z15 <= 16'd48;
		81: z15 <= 16'd41;
		82: z15 <= -16'd92;
		83: z15 <= -16'd128;
		84: z15 <= 16'd127;
		85: z15 <= 16'd45;
		86: z15 <= 16'd93;
		87: z15 <= 16'd2;
		88: z15 <= 16'd15;
		89: z15 <= 16'd5;
		90: z15 <= -16'd85;
		91: z15 <= 16'd41;
		92: z15 <= 16'd107;
		93: z15 <= 16'd68;
		94: z15 <= 16'd113;
		95: z15 <= 16'd55;
		96: z15 <= -16'd48;
		97: z15 <= -16'd82;
		98: z15 <= -16'd50;
		99: z15 <= 16'd94;
		100: z15 <= 16'd10;
		101: z15 <= 16'd55;
		102: z15 <= -16'd40;
		103: z15 <= -16'd20;
		104: z15 <= 16'd102;
		105: z15 <= 16'd22;
		106: z15 <= 16'd47;
		107: z15 <= -16'd12;
		108: z15 <= -16'd39;
		109: z15 <= -16'd21;
		110: z15 <= -16'd85;
		111: z15 <= -16'd118;
		112: z15 <= -16'd108;
		113: z15 <= -16'd48;
		114: z15 <= -16'd118;
		115: z15 <= -16'd109;
		116: z15 <= 16'd125;
		117: z15 <= 16'd103;
		118: z15 <= 16'd21;
		119: z15 <= 16'd12;
		120: z15 <= -16'd19;
		121: z15 <= 16'd64;
		122: z15 <= -16'd75;
		123: z15 <= -16'd40;
		124: z15 <= 16'd4;
		125: z15 <= -16'd89;
		126: z15 <= -16'd113;
		127: z15 <= 16'd85;
		endcase
	end
endmodule

