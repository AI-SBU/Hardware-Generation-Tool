module fc_16_12_20_0_1(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 16;
	parameter N = 12;
	parameter T = 20;
	parameter R = 0;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned[7 : 0] addr_w;
	logic unsigned[3 : 0] addr_x;
	logic signed [19 : 0] v_out, m_out;
	logic unsigned wr_en_x;
	logic unsigned clear_acc;
	logic unsigned en_acc;

	controlFSM #(16,12) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr_w), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid));

	datapath #(20, 0) datapathMod(.clk(clk), .reset(reset), .m_out(m_out), .v_out(v_out),
									.en_acc(en_acc), .output_data(output_data), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	memory #(20, 12 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	fc_16_12_20_0_1_W_rom  matrixRom(.clk(clk), .addr(addr_w), .z(m_out));

endmodule

module fc_16_12_20_0_1_W_rom(clk, addr, z);
   input clk;
   input [7:0] addr;
   output logic signed [19:0] z;
   always_ff @(posedge clk) begin
      case(addr)
        0: z <= 20'd216;
        1: z <= 20'd116;
        2: z <= 20'd128;
        3: z <= 20'd38;
        4: z <= -20'd263;
        5: z <= 20'd470;
        6: z <= -20'd412;
        7: z <= 20'd367;
        8: z <= -20'd114;
        9: z <= 20'd458;
        10: z <= -20'd66;
        11: z <= -20'd86;
        12: z <= -20'd163;
        13: z <= -20'd150;
        14: z <= 20'd179;
        15: z <= -20'd459;
        16: z <= 20'd67;
        17: z <= -20'd51;
        18: z <= -20'd24;
        19: z <= -20'd442;
        20: z <= 20'd467;
        21: z <= -20'd81;
        22: z <= -20'd17;
        23: z <= 20'd141;
        24: z <= -20'd163;
        25: z <= -20'd293;
        26: z <= -20'd281;
        27: z <= 20'd34;
        28: z <= 20'd250;
        29: z <= 20'd102;
        30: z <= 20'd510;
        31: z <= -20'd45;
        32: z <= -20'd293;
        33: z <= 20'd126;
        34: z <= 20'd505;
        35: z <= -20'd44;
        36: z <= 20'd84;
        37: z <= -20'd419;
        38: z <= -20'd189;
        39: z <= 20'd482;
        40: z <= -20'd472;
        41: z <= 20'd258;
        42: z <= -20'd116;
        43: z <= -20'd123;
        44: z <= -20'd404;
        45: z <= -20'd448;
        46: z <= -20'd70;
        47: z <= 20'd175;
        48: z <= 20'd13;
        49: z <= 20'd419;
        50: z <= 20'd245;
        51: z <= -20'd32;
        52: z <= -20'd174;
        53: z <= -20'd283;
        54: z <= -20'd403;
        55: z <= 20'd175;
        56: z <= -20'd64;
        57: z <= -20'd172;
        58: z <= -20'd303;
        59: z <= -20'd326;
        60: z <= 20'd443;
        61: z <= -20'd305;
        62: z <= 20'd141;
        63: z <= -20'd362;
        64: z <= 20'd333;
        65: z <= 20'd134;
        66: z <= 20'd106;
        67: z <= -20'd94;
        68: z <= 20'd228;
        69: z <= 20'd430;
        70: z <= -20'd124;
        71: z <= 20'd268;
        72: z <= 20'd176;
        73: z <= 20'd273;
        74: z <= -20'd367;
        75: z <= 20'd284;
        76: z <= 20'd337;
        77: z <= 20'd76;
        78: z <= -20'd53;
        79: z <= -20'd162;
        80: z <= -20'd17;
        81: z <= -20'd320;
        82: z <= 20'd318;
        83: z <= 20'd321;
        84: z <= -20'd91;
        85: z <= 20'd427;
        86: z <= -20'd16;
        87: z <= 20'd357;
        88: z <= -20'd256;
        89: z <= 20'd194;
        90: z <= -20'd480;
        91: z <= -20'd325;
        92: z <= 20'd401;
        93: z <= 20'd173;
        94: z <= -20'd175;
        95: z <= 20'd223;
        96: z <= -20'd204;
        97: z <= 20'd443;
        98: z <= -20'd383;
        99: z <= -20'd488;
        100: z <= 20'd361;
        101: z <= 20'd5;
        102: z <= 20'd292;
        103: z <= 20'd25;
        104: z <= -20'd234;
        105: z <= 20'd437;
        106: z <= -20'd203;
        107: z <= -20'd409;
        108: z <= 20'd1;
        109: z <= 20'd256;
        110: z <= -20'd59;
        111: z <= 20'd496;
        112: z <= 20'd449;
        113: z <= -20'd253;
        114: z <= 20'd305;
        115: z <= -20'd154;
        116: z <= -20'd337;
        117: z <= -20'd222;
        118: z <= -20'd308;
        119: z <= -20'd81;
        120: z <= 20'd484;
        121: z <= -20'd276;
        122: z <= 20'd106;
        123: z <= 20'd373;
        124: z <= 20'd409;
        125: z <= 20'd443;
        126: z <= 20'd84;
        127: z <= -20'd307;
        128: z <= 20'd374;
        129: z <= 20'd213;
        130: z <= -20'd283;
        131: z <= 20'd224;
        132: z <= -20'd293;
        133: z <= -20'd503;
        134: z <= -20'd263;
        135: z <= -20'd15;
        136: z <= 20'd447;
        137: z <= 20'd47;
        138: z <= 20'd89;
        139: z <= -20'd64;
        140: z <= -20'd209;
        141: z <= -20'd482;
        142: z <= -20'd79;
        143: z <= -20'd272;
        144: z <= -20'd222;
        145: z <= -20'd286;
        146: z <= 20'd87;
        147: z <= -20'd47;
        148: z <= 20'd4;
        149: z <= 20'd291;
        150: z <= 20'd384;
        151: z <= -20'd24;
        152: z <= -20'd497;
        153: z <= -20'd22;
        154: z <= -20'd162;
        155: z <= 20'd424;
        156: z <= -20'd91;
        157: z <= 20'd434;
        158: z <= -20'd394;
        159: z <= -20'd229;
        160: z <= 20'd136;
        161: z <= -20'd165;
        162: z <= 20'd507;
        163: z <= 20'd355;
        164: z <= -20'd155;
        165: z <= -20'd267;
        166: z <= -20'd172;
        167: z <= -20'd220;
        168: z <= 20'd292;
        169: z <= 20'd429;
        170: z <= 20'd228;
        171: z <= -20'd429;
        172: z <= 20'd460;
        173: z <= -20'd363;
        174: z <= -20'd188;
        175: z <= -20'd274;
        176: z <= -20'd136;
        177: z <= 20'd411;
        178: z <= 20'd191;
        179: z <= 20'd380;
        180: z <= 20'd190;
        181: z <= 20'd63;
        182: z <= -20'd155;
        183: z <= 20'd205;
        184: z <= -20'd471;
        185: z <= 20'd195;
        186: z <= 20'd117;
        187: z <= -20'd50;
        188: z <= 20'd117;
        189: z <= 20'd235;
        190: z <= 20'd233;
        191: z <= -20'd259;
      endcase
   end
endmodule

