`include "controlFSM.sv"
`include "datapath.sv"
`include "memory.sv"

module fc_16_8_16_1_8(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 16;
	parameter N = 8;
	parameter T = 16;
	parameter R = 1;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned [2 : 0] sel;

	logic signed [T-1 : 0] parallel_out0;
	logic signed [T-1 : 0] parallel_out1;
	logic signed [T-1 : 0] parallel_out2;
	logic signed [T-1 : 0] parallel_out3;
	logic signed [T-1 : 0] parallel_out4;
	logic signed [T-1 : 0] parallel_out5;
	logic signed [T-1 : 0] parallel_out6;
	logic signed [T-1 : 0] parallel_out7;

	logic unsigned[2 : 0] addr_x;
	logic signed [15 : 0] v_out;
	logic unsigned wr_en_x;

	logic unsigned[6 : 0] addr;

	logic unsigned[6 : 0] addr_w0;
	logic signed [15 : 0] m_out0;

	logic unsigned[6 : 0] addr_w1;
	logic signed [15 : 0] m_out1;

	logic unsigned[6 : 0] addr_w2;
	logic signed [15 : 0] m_out2;

	logic unsigned[6 : 0] addr_w3;
	logic signed [15 : 0] m_out3;

	logic unsigned[6 : 0] addr_w4;
	logic signed [15 : 0] m_out4;

	logic unsigned[6 : 0] addr_w5;
	logic signed [15 : 0] m_out5;

	logic unsigned[6 : 0] addr_w6;
	logic signed [15 : 0] m_out6;

	logic unsigned[6 : 0] addr_w7;
	logic signed [15 : 0] m_out7;

	logic unsigned clear_acc;
	logic unsigned en_acc;

	always_comb begin
		addr_w0 = addr + 0;
		addr_w1 = addr + 8;
		addr_w2 = addr + 16;
		addr_w3 = addr + 24;
		addr_w4 = addr + 32;
		addr_w5 = addr + 40;
		addr_w6 = addr + 48;
		addr_w7 = addr + 56;
	end

	controlFSM #(16,8,8) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid), .countToP(sel));

	memory #(16, 8 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	mux #(16, 8) muxMod(.parallel_out0(parallel_out0), .parallel_out1(parallel_out1), .parallel_out2(parallel_out2), .parallel_out3(parallel_out3), .parallel_out4(parallel_out4), .parallel_out5(parallel_out5), .parallel_out6(parallel_out6), .parallel_out7(parallel_out7), .sel(sel), .f(output_data));

	datapath #(16, 1) datapathMod0(.clk(clk), .reset(reset), .m_out(m_out0), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out0), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod1(.clk(clk), .reset(reset), .m_out(m_out1), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out1), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod2(.clk(clk), .reset(reset), .m_out(m_out2), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out2), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod3(.clk(clk), .reset(reset), .m_out(m_out3), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out3), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod4(.clk(clk), .reset(reset), .m_out(m_out4), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out4), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod5(.clk(clk), .reset(reset), .m_out(m_out5), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out5), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod6(.clk(clk), .reset(reset), .m_out(m_out6), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out6), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod7(.clk(clk), .reset(reset), .m_out(m_out7), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out7), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	fc_16_8_16_1_8_W_rom  matrixRom(.clk(clk),.addr0(addr_w0), .addr1(addr_w1), .addr2(addr_w2), .addr3(addr_w3), .addr4(addr_w4), .addr5(addr_w5), .addr6(addr_w6), .addr7(addr_w7), .z0(m_out0), .z1(m_out1), .z2(m_out2), .z3(m_out3), .z4(m_out4), .z5(m_out5), .z6(m_out6), .z7(m_out7));

endmodule

module mux(parallel_out0, parallel_out1, parallel_out2, parallel_out3, parallel_out4, parallel_out5, parallel_out6, parallel_out7, sel, f);
	parameter T = 16;
	parameter P = 8;

	output signed [T-1 : 0] f;
	input logic unsigned [2 : 0] sel;
	input signed [T-1 : 0] parallel_out0;
	input signed [T-1 : 0] parallel_out1;
	input signed [T-1 : 0] parallel_out2;
	input signed [T-1 : 0] parallel_out3;
	input signed [T-1 : 0] parallel_out4;
	input signed [T-1 : 0] parallel_out5;
	input signed [T-1 : 0] parallel_out6;
	input signed [T-1 : 0] parallel_out7;
	logic unsigned [P*T-1 : 0] array;
	assign  array = {parallel_out0[15 : 0], parallel_out1[15 : 0], parallel_out2[15 : 0], parallel_out3[15 : 0], parallel_out4[15 : 0], parallel_out5[15 : 0], parallel_out6[15 : 0], parallel_out7[15: 0]};

	assign f = (sel == 0) ? parallel_out0 : 
			(sel == 1) ? parallel_out1 : 
			(sel == 2) ? parallel_out2 : 
			(sel == 3) ? parallel_out3 : 
			(sel == 4) ? parallel_out4 : 
			(sel == 5) ? parallel_out5 : 
			(sel == 6) ? parallel_out6 : 
			(sel == 7) ? parallel_out7 : 16'bz;
endmodule

module fc_16_8_16_1_8_W_rom(clk, addr0, addr1, addr2, addr3, addr4, addr5, addr6, addr7, z0, z1, z2, z3, z4, z5, z6, z7);
	input clk;
	input [6:0] addr0;
	input [6:0] addr1;
	input [6:0] addr2;
	input [6:0] addr3;
	input [6:0] addr4;
	input [6:0] addr5;
	input [6:0] addr6;
	input [6:0] addr7;
	output logic signed [15:0] z0;
	output logic signed [15:0] z1;
	output logic signed [15:0] z2;
	output logic signed [15:0] z3;
	output logic signed [15:0] z4;
	output logic signed [15:0] z5;
	output logic signed [15:0] z6;
	output logic signed [15:0] z7;
	always_ff @(posedge clk) begin
		case(addr0)
		0: z0 <= 16'd119;
		1: z0 <= 16'd104;
		2: z0 <= -16'd111;
		3: z0 <= 16'd114;
		4: z0 <= -16'd1;
		5: z0 <= -16'd6;
		6: z0 <= 16'd39;
		7: z0 <= -16'd91;
		8: z0 <= -16'd21;
		9: z0 <= -16'd60;
		10: z0 <= -16'd57;
		11: z0 <= 16'd28;
		12: z0 <= 16'd21;
		13: z0 <= -16'd55;
		14: z0 <= -16'd26;
		15: z0 <= 16'd77;
		16: z0 <= 16'd17;
		17: z0 <= -16'd39;
		18: z0 <= -16'd3;
		19: z0 <= -16'd92;
		20: z0 <= -16'd79;
		21: z0 <= 16'd123;
		22: z0 <= 16'd59;
		23: z0 <= 16'd83;
		24: z0 <= -16'd28;
		25: z0 <= 16'd74;
		26: z0 <= 16'd67;
		27: z0 <= 16'd21;
		28: z0 <= -16'd109;
		29: z0 <= -16'd18;
		30: z0 <= -16'd30;
		31: z0 <= -16'd118;
		32: z0 <= -16'd42;
		33: z0 <= -16'd13;
		34: z0 <= 16'd124;
		35: z0 <= 16'd85;
		36: z0 <= 16'd109;
		37: z0 <= 16'd36;
		38: z0 <= 16'd122;
		39: z0 <= -16'd39;
		40: z0 <= 16'd104;
		41: z0 <= -16'd62;
		42: z0 <= 16'd117;
		43: z0 <= -16'd3;
		44: z0 <= 16'd11;
		45: z0 <= -16'd36;
		46: z0 <= -16'd54;
		47: z0 <= -16'd100;
		48: z0 <= 16'd53;
		49: z0 <= 16'd71;
		50: z0 <= -16'd63;
		51: z0 <= 16'd102;
		52: z0 <= 16'd67;
		53: z0 <= 16'd124;
		54: z0 <= 16'd58;
		55: z0 <= -16'd89;
		56: z0 <= 16'd70;
		57: z0 <= -16'd3;
		58: z0 <= 16'd61;
		59: z0 <= 16'd89;
		60: z0 <= 16'd108;
		61: z0 <= -16'd97;
		62: z0 <= 16'd100;
		63: z0 <= -16'd62;
		64: z0 <= 16'd18;
		65: z0 <= 16'd96;
		66: z0 <= -16'd104;
		67: z0 <= 16'd0;
		68: z0 <= 16'd4;
		69: z0 <= -16'd110;
		70: z0 <= 16'd89;
		71: z0 <= -16'd20;
		72: z0 <= -16'd44;
		73: z0 <= 16'd78;
		74: z0 <= 16'd106;
		75: z0 <= 16'd96;
		76: z0 <= -16'd86;
		77: z0 <= -16'd76;
		78: z0 <= 16'd124;
		79: z0 <= 16'd96;
		80: z0 <= 16'd124;
		81: z0 <= -16'd67;
		82: z0 <= 16'd70;
		83: z0 <= 16'd63;
		84: z0 <= -16'd71;
		85: z0 <= 16'd0;
		86: z0 <= 16'd102;
		87: z0 <= 16'd127;
		88: z0 <= 16'd126;
		89: z0 <= 16'd35;
		90: z0 <= 16'd89;
		91: z0 <= 16'd106;
		92: z0 <= 16'd66;
		93: z0 <= 16'd61;
		94: z0 <= -16'd84;
		95: z0 <= -16'd43;
		96: z0 <= 16'd29;
		97: z0 <= -16'd60;
		98: z0 <= 16'd85;
		99: z0 <= -16'd94;
		100: z0 <= -16'd41;
		101: z0 <= 16'd46;
		102: z0 <= 16'd14;
		103: z0 <= 16'd43;
		104: z0 <= -16'd4;
		105: z0 <= -16'd8;
		106: z0 <= 16'd11;
		107: z0 <= 16'd39;
		108: z0 <= 16'd45;
		109: z0 <= 16'd8;
		110: z0 <= 16'd7;
		111: z0 <= 16'd41;
		112: z0 <= 16'd69;
		113: z0 <= -16'd51;
		114: z0 <= -16'd24;
		115: z0 <= 16'd127;
		116: z0 <= 16'd78;
		117: z0 <= -16'd50;
		118: z0 <= 16'd126;
		119: z0 <= 16'd76;
		120: z0 <= 16'd114;
		121: z0 <= 16'd87;
		122: z0 <= 16'd54;
		123: z0 <= 16'd52;
		124: z0 <= 16'd20;
		125: z0 <= 16'd98;
		126: z0 <= -16'd119;
		127: z0 <= -16'd78;
		endcase
		case(addr1)
		0: z1 <= 16'd119;
		1: z1 <= 16'd104;
		2: z1 <= -16'd111;
		3: z1 <= 16'd114;
		4: z1 <= -16'd1;
		5: z1 <= -16'd6;
		6: z1 <= 16'd39;
		7: z1 <= -16'd91;
		8: z1 <= -16'd21;
		9: z1 <= -16'd60;
		10: z1 <= -16'd57;
		11: z1 <= 16'd28;
		12: z1 <= 16'd21;
		13: z1 <= -16'd55;
		14: z1 <= -16'd26;
		15: z1 <= 16'd77;
		16: z1 <= 16'd17;
		17: z1 <= -16'd39;
		18: z1 <= -16'd3;
		19: z1 <= -16'd92;
		20: z1 <= -16'd79;
		21: z1 <= 16'd123;
		22: z1 <= 16'd59;
		23: z1 <= 16'd83;
		24: z1 <= -16'd28;
		25: z1 <= 16'd74;
		26: z1 <= 16'd67;
		27: z1 <= 16'd21;
		28: z1 <= -16'd109;
		29: z1 <= -16'd18;
		30: z1 <= -16'd30;
		31: z1 <= -16'd118;
		32: z1 <= -16'd42;
		33: z1 <= -16'd13;
		34: z1 <= 16'd124;
		35: z1 <= 16'd85;
		36: z1 <= 16'd109;
		37: z1 <= 16'd36;
		38: z1 <= 16'd122;
		39: z1 <= -16'd39;
		40: z1 <= 16'd104;
		41: z1 <= -16'd62;
		42: z1 <= 16'd117;
		43: z1 <= -16'd3;
		44: z1 <= 16'd11;
		45: z1 <= -16'd36;
		46: z1 <= -16'd54;
		47: z1 <= -16'd100;
		48: z1 <= 16'd53;
		49: z1 <= 16'd71;
		50: z1 <= -16'd63;
		51: z1 <= 16'd102;
		52: z1 <= 16'd67;
		53: z1 <= 16'd124;
		54: z1 <= 16'd58;
		55: z1 <= -16'd89;
		56: z1 <= 16'd70;
		57: z1 <= -16'd3;
		58: z1 <= 16'd61;
		59: z1 <= 16'd89;
		60: z1 <= 16'd108;
		61: z1 <= -16'd97;
		62: z1 <= 16'd100;
		63: z1 <= -16'd62;
		64: z1 <= 16'd18;
		65: z1 <= 16'd96;
		66: z1 <= -16'd104;
		67: z1 <= 16'd0;
		68: z1 <= 16'd4;
		69: z1 <= -16'd110;
		70: z1 <= 16'd89;
		71: z1 <= -16'd20;
		72: z1 <= -16'd44;
		73: z1 <= 16'd78;
		74: z1 <= 16'd106;
		75: z1 <= 16'd96;
		76: z1 <= -16'd86;
		77: z1 <= -16'd76;
		78: z1 <= 16'd124;
		79: z1 <= 16'd96;
		80: z1 <= 16'd124;
		81: z1 <= -16'd67;
		82: z1 <= 16'd70;
		83: z1 <= 16'd63;
		84: z1 <= -16'd71;
		85: z1 <= 16'd0;
		86: z1 <= 16'd102;
		87: z1 <= 16'd127;
		88: z1 <= 16'd126;
		89: z1 <= 16'd35;
		90: z1 <= 16'd89;
		91: z1 <= 16'd106;
		92: z1 <= 16'd66;
		93: z1 <= 16'd61;
		94: z1 <= -16'd84;
		95: z1 <= -16'd43;
		96: z1 <= 16'd29;
		97: z1 <= -16'd60;
		98: z1 <= 16'd85;
		99: z1 <= -16'd94;
		100: z1 <= -16'd41;
		101: z1 <= 16'd46;
		102: z1 <= 16'd14;
		103: z1 <= 16'd43;
		104: z1 <= -16'd4;
		105: z1 <= -16'd8;
		106: z1 <= 16'd11;
		107: z1 <= 16'd39;
		108: z1 <= 16'd45;
		109: z1 <= 16'd8;
		110: z1 <= 16'd7;
		111: z1 <= 16'd41;
		112: z1 <= 16'd69;
		113: z1 <= -16'd51;
		114: z1 <= -16'd24;
		115: z1 <= 16'd127;
		116: z1 <= 16'd78;
		117: z1 <= -16'd50;
		118: z1 <= 16'd126;
		119: z1 <= 16'd76;
		120: z1 <= 16'd114;
		121: z1 <= 16'd87;
		122: z1 <= 16'd54;
		123: z1 <= 16'd52;
		124: z1 <= 16'd20;
		125: z1 <= 16'd98;
		126: z1 <= -16'd119;
		127: z1 <= -16'd78;
		endcase
		case(addr2)
		0: z2 <= 16'd119;
		1: z2 <= 16'd104;
		2: z2 <= -16'd111;
		3: z2 <= 16'd114;
		4: z2 <= -16'd1;
		5: z2 <= -16'd6;
		6: z2 <= 16'd39;
		7: z2 <= -16'd91;
		8: z2 <= -16'd21;
		9: z2 <= -16'd60;
		10: z2 <= -16'd57;
		11: z2 <= 16'd28;
		12: z2 <= 16'd21;
		13: z2 <= -16'd55;
		14: z2 <= -16'd26;
		15: z2 <= 16'd77;
		16: z2 <= 16'd17;
		17: z2 <= -16'd39;
		18: z2 <= -16'd3;
		19: z2 <= -16'd92;
		20: z2 <= -16'd79;
		21: z2 <= 16'd123;
		22: z2 <= 16'd59;
		23: z2 <= 16'd83;
		24: z2 <= -16'd28;
		25: z2 <= 16'd74;
		26: z2 <= 16'd67;
		27: z2 <= 16'd21;
		28: z2 <= -16'd109;
		29: z2 <= -16'd18;
		30: z2 <= -16'd30;
		31: z2 <= -16'd118;
		32: z2 <= -16'd42;
		33: z2 <= -16'd13;
		34: z2 <= 16'd124;
		35: z2 <= 16'd85;
		36: z2 <= 16'd109;
		37: z2 <= 16'd36;
		38: z2 <= 16'd122;
		39: z2 <= -16'd39;
		40: z2 <= 16'd104;
		41: z2 <= -16'd62;
		42: z2 <= 16'd117;
		43: z2 <= -16'd3;
		44: z2 <= 16'd11;
		45: z2 <= -16'd36;
		46: z2 <= -16'd54;
		47: z2 <= -16'd100;
		48: z2 <= 16'd53;
		49: z2 <= 16'd71;
		50: z2 <= -16'd63;
		51: z2 <= 16'd102;
		52: z2 <= 16'd67;
		53: z2 <= 16'd124;
		54: z2 <= 16'd58;
		55: z2 <= -16'd89;
		56: z2 <= 16'd70;
		57: z2 <= -16'd3;
		58: z2 <= 16'd61;
		59: z2 <= 16'd89;
		60: z2 <= 16'd108;
		61: z2 <= -16'd97;
		62: z2 <= 16'd100;
		63: z2 <= -16'd62;
		64: z2 <= 16'd18;
		65: z2 <= 16'd96;
		66: z2 <= -16'd104;
		67: z2 <= 16'd0;
		68: z2 <= 16'd4;
		69: z2 <= -16'd110;
		70: z2 <= 16'd89;
		71: z2 <= -16'd20;
		72: z2 <= -16'd44;
		73: z2 <= 16'd78;
		74: z2 <= 16'd106;
		75: z2 <= 16'd96;
		76: z2 <= -16'd86;
		77: z2 <= -16'd76;
		78: z2 <= 16'd124;
		79: z2 <= 16'd96;
		80: z2 <= 16'd124;
		81: z2 <= -16'd67;
		82: z2 <= 16'd70;
		83: z2 <= 16'd63;
		84: z2 <= -16'd71;
		85: z2 <= 16'd0;
		86: z2 <= 16'd102;
		87: z2 <= 16'd127;
		88: z2 <= 16'd126;
		89: z2 <= 16'd35;
		90: z2 <= 16'd89;
		91: z2 <= 16'd106;
		92: z2 <= 16'd66;
		93: z2 <= 16'd61;
		94: z2 <= -16'd84;
		95: z2 <= -16'd43;
		96: z2 <= 16'd29;
		97: z2 <= -16'd60;
		98: z2 <= 16'd85;
		99: z2 <= -16'd94;
		100: z2 <= -16'd41;
		101: z2 <= 16'd46;
		102: z2 <= 16'd14;
		103: z2 <= 16'd43;
		104: z2 <= -16'd4;
		105: z2 <= -16'd8;
		106: z2 <= 16'd11;
		107: z2 <= 16'd39;
		108: z2 <= 16'd45;
		109: z2 <= 16'd8;
		110: z2 <= 16'd7;
		111: z2 <= 16'd41;
		112: z2 <= 16'd69;
		113: z2 <= -16'd51;
		114: z2 <= -16'd24;
		115: z2 <= 16'd127;
		116: z2 <= 16'd78;
		117: z2 <= -16'd50;
		118: z2 <= 16'd126;
		119: z2 <= 16'd76;
		120: z2 <= 16'd114;
		121: z2 <= 16'd87;
		122: z2 <= 16'd54;
		123: z2 <= 16'd52;
		124: z2 <= 16'd20;
		125: z2 <= 16'd98;
		126: z2 <= -16'd119;
		127: z2 <= -16'd78;
		endcase
		case(addr3)
		0: z3 <= 16'd119;
		1: z3 <= 16'd104;
		2: z3 <= -16'd111;
		3: z3 <= 16'd114;
		4: z3 <= -16'd1;
		5: z3 <= -16'd6;
		6: z3 <= 16'd39;
		7: z3 <= -16'd91;
		8: z3 <= -16'd21;
		9: z3 <= -16'd60;
		10: z3 <= -16'd57;
		11: z3 <= 16'd28;
		12: z3 <= 16'd21;
		13: z3 <= -16'd55;
		14: z3 <= -16'd26;
		15: z3 <= 16'd77;
		16: z3 <= 16'd17;
		17: z3 <= -16'd39;
		18: z3 <= -16'd3;
		19: z3 <= -16'd92;
		20: z3 <= -16'd79;
		21: z3 <= 16'd123;
		22: z3 <= 16'd59;
		23: z3 <= 16'd83;
		24: z3 <= -16'd28;
		25: z3 <= 16'd74;
		26: z3 <= 16'd67;
		27: z3 <= 16'd21;
		28: z3 <= -16'd109;
		29: z3 <= -16'd18;
		30: z3 <= -16'd30;
		31: z3 <= -16'd118;
		32: z3 <= -16'd42;
		33: z3 <= -16'd13;
		34: z3 <= 16'd124;
		35: z3 <= 16'd85;
		36: z3 <= 16'd109;
		37: z3 <= 16'd36;
		38: z3 <= 16'd122;
		39: z3 <= -16'd39;
		40: z3 <= 16'd104;
		41: z3 <= -16'd62;
		42: z3 <= 16'd117;
		43: z3 <= -16'd3;
		44: z3 <= 16'd11;
		45: z3 <= -16'd36;
		46: z3 <= -16'd54;
		47: z3 <= -16'd100;
		48: z3 <= 16'd53;
		49: z3 <= 16'd71;
		50: z3 <= -16'd63;
		51: z3 <= 16'd102;
		52: z3 <= 16'd67;
		53: z3 <= 16'd124;
		54: z3 <= 16'd58;
		55: z3 <= -16'd89;
		56: z3 <= 16'd70;
		57: z3 <= -16'd3;
		58: z3 <= 16'd61;
		59: z3 <= 16'd89;
		60: z3 <= 16'd108;
		61: z3 <= -16'd97;
		62: z3 <= 16'd100;
		63: z3 <= -16'd62;
		64: z3 <= 16'd18;
		65: z3 <= 16'd96;
		66: z3 <= -16'd104;
		67: z3 <= 16'd0;
		68: z3 <= 16'd4;
		69: z3 <= -16'd110;
		70: z3 <= 16'd89;
		71: z3 <= -16'd20;
		72: z3 <= -16'd44;
		73: z3 <= 16'd78;
		74: z3 <= 16'd106;
		75: z3 <= 16'd96;
		76: z3 <= -16'd86;
		77: z3 <= -16'd76;
		78: z3 <= 16'd124;
		79: z3 <= 16'd96;
		80: z3 <= 16'd124;
		81: z3 <= -16'd67;
		82: z3 <= 16'd70;
		83: z3 <= 16'd63;
		84: z3 <= -16'd71;
		85: z3 <= 16'd0;
		86: z3 <= 16'd102;
		87: z3 <= 16'd127;
		88: z3 <= 16'd126;
		89: z3 <= 16'd35;
		90: z3 <= 16'd89;
		91: z3 <= 16'd106;
		92: z3 <= 16'd66;
		93: z3 <= 16'd61;
		94: z3 <= -16'd84;
		95: z3 <= -16'd43;
		96: z3 <= 16'd29;
		97: z3 <= -16'd60;
		98: z3 <= 16'd85;
		99: z3 <= -16'd94;
		100: z3 <= -16'd41;
		101: z3 <= 16'd46;
		102: z3 <= 16'd14;
		103: z3 <= 16'd43;
		104: z3 <= -16'd4;
		105: z3 <= -16'd8;
		106: z3 <= 16'd11;
		107: z3 <= 16'd39;
		108: z3 <= 16'd45;
		109: z3 <= 16'd8;
		110: z3 <= 16'd7;
		111: z3 <= 16'd41;
		112: z3 <= 16'd69;
		113: z3 <= -16'd51;
		114: z3 <= -16'd24;
		115: z3 <= 16'd127;
		116: z3 <= 16'd78;
		117: z3 <= -16'd50;
		118: z3 <= 16'd126;
		119: z3 <= 16'd76;
		120: z3 <= 16'd114;
		121: z3 <= 16'd87;
		122: z3 <= 16'd54;
		123: z3 <= 16'd52;
		124: z3 <= 16'd20;
		125: z3 <= 16'd98;
		126: z3 <= -16'd119;
		127: z3 <= -16'd78;
		endcase
		case(addr4)
		0: z4 <= 16'd119;
		1: z4 <= 16'd104;
		2: z4 <= -16'd111;
		3: z4 <= 16'd114;
		4: z4 <= -16'd1;
		5: z4 <= -16'd6;
		6: z4 <= 16'd39;
		7: z4 <= -16'd91;
		8: z4 <= -16'd21;
		9: z4 <= -16'd60;
		10: z4 <= -16'd57;
		11: z4 <= 16'd28;
		12: z4 <= 16'd21;
		13: z4 <= -16'd55;
		14: z4 <= -16'd26;
		15: z4 <= 16'd77;
		16: z4 <= 16'd17;
		17: z4 <= -16'd39;
		18: z4 <= -16'd3;
		19: z4 <= -16'd92;
		20: z4 <= -16'd79;
		21: z4 <= 16'd123;
		22: z4 <= 16'd59;
		23: z4 <= 16'd83;
		24: z4 <= -16'd28;
		25: z4 <= 16'd74;
		26: z4 <= 16'd67;
		27: z4 <= 16'd21;
		28: z4 <= -16'd109;
		29: z4 <= -16'd18;
		30: z4 <= -16'd30;
		31: z4 <= -16'd118;
		32: z4 <= -16'd42;
		33: z4 <= -16'd13;
		34: z4 <= 16'd124;
		35: z4 <= 16'd85;
		36: z4 <= 16'd109;
		37: z4 <= 16'd36;
		38: z4 <= 16'd122;
		39: z4 <= -16'd39;
		40: z4 <= 16'd104;
		41: z4 <= -16'd62;
		42: z4 <= 16'd117;
		43: z4 <= -16'd3;
		44: z4 <= 16'd11;
		45: z4 <= -16'd36;
		46: z4 <= -16'd54;
		47: z4 <= -16'd100;
		48: z4 <= 16'd53;
		49: z4 <= 16'd71;
		50: z4 <= -16'd63;
		51: z4 <= 16'd102;
		52: z4 <= 16'd67;
		53: z4 <= 16'd124;
		54: z4 <= 16'd58;
		55: z4 <= -16'd89;
		56: z4 <= 16'd70;
		57: z4 <= -16'd3;
		58: z4 <= 16'd61;
		59: z4 <= 16'd89;
		60: z4 <= 16'd108;
		61: z4 <= -16'd97;
		62: z4 <= 16'd100;
		63: z4 <= -16'd62;
		64: z4 <= 16'd18;
		65: z4 <= 16'd96;
		66: z4 <= -16'd104;
		67: z4 <= 16'd0;
		68: z4 <= 16'd4;
		69: z4 <= -16'd110;
		70: z4 <= 16'd89;
		71: z4 <= -16'd20;
		72: z4 <= -16'd44;
		73: z4 <= 16'd78;
		74: z4 <= 16'd106;
		75: z4 <= 16'd96;
		76: z4 <= -16'd86;
		77: z4 <= -16'd76;
		78: z4 <= 16'd124;
		79: z4 <= 16'd96;
		80: z4 <= 16'd124;
		81: z4 <= -16'd67;
		82: z4 <= 16'd70;
		83: z4 <= 16'd63;
		84: z4 <= -16'd71;
		85: z4 <= 16'd0;
		86: z4 <= 16'd102;
		87: z4 <= 16'd127;
		88: z4 <= 16'd126;
		89: z4 <= 16'd35;
		90: z4 <= 16'd89;
		91: z4 <= 16'd106;
		92: z4 <= 16'd66;
		93: z4 <= 16'd61;
		94: z4 <= -16'd84;
		95: z4 <= -16'd43;
		96: z4 <= 16'd29;
		97: z4 <= -16'd60;
		98: z4 <= 16'd85;
		99: z4 <= -16'd94;
		100: z4 <= -16'd41;
		101: z4 <= 16'd46;
		102: z4 <= 16'd14;
		103: z4 <= 16'd43;
		104: z4 <= -16'd4;
		105: z4 <= -16'd8;
		106: z4 <= 16'd11;
		107: z4 <= 16'd39;
		108: z4 <= 16'd45;
		109: z4 <= 16'd8;
		110: z4 <= 16'd7;
		111: z4 <= 16'd41;
		112: z4 <= 16'd69;
		113: z4 <= -16'd51;
		114: z4 <= -16'd24;
		115: z4 <= 16'd127;
		116: z4 <= 16'd78;
		117: z4 <= -16'd50;
		118: z4 <= 16'd126;
		119: z4 <= 16'd76;
		120: z4 <= 16'd114;
		121: z4 <= 16'd87;
		122: z4 <= 16'd54;
		123: z4 <= 16'd52;
		124: z4 <= 16'd20;
		125: z4 <= 16'd98;
		126: z4 <= -16'd119;
		127: z4 <= -16'd78;
		endcase
		case(addr5)
		0: z5 <= 16'd119;
		1: z5 <= 16'd104;
		2: z5 <= -16'd111;
		3: z5 <= 16'd114;
		4: z5 <= -16'd1;
		5: z5 <= -16'd6;
		6: z5 <= 16'd39;
		7: z5 <= -16'd91;
		8: z5 <= -16'd21;
		9: z5 <= -16'd60;
		10: z5 <= -16'd57;
		11: z5 <= 16'd28;
		12: z5 <= 16'd21;
		13: z5 <= -16'd55;
		14: z5 <= -16'd26;
		15: z5 <= 16'd77;
		16: z5 <= 16'd17;
		17: z5 <= -16'd39;
		18: z5 <= -16'd3;
		19: z5 <= -16'd92;
		20: z5 <= -16'd79;
		21: z5 <= 16'd123;
		22: z5 <= 16'd59;
		23: z5 <= 16'd83;
		24: z5 <= -16'd28;
		25: z5 <= 16'd74;
		26: z5 <= 16'd67;
		27: z5 <= 16'd21;
		28: z5 <= -16'd109;
		29: z5 <= -16'd18;
		30: z5 <= -16'd30;
		31: z5 <= -16'd118;
		32: z5 <= -16'd42;
		33: z5 <= -16'd13;
		34: z5 <= 16'd124;
		35: z5 <= 16'd85;
		36: z5 <= 16'd109;
		37: z5 <= 16'd36;
		38: z5 <= 16'd122;
		39: z5 <= -16'd39;
		40: z5 <= 16'd104;
		41: z5 <= -16'd62;
		42: z5 <= 16'd117;
		43: z5 <= -16'd3;
		44: z5 <= 16'd11;
		45: z5 <= -16'd36;
		46: z5 <= -16'd54;
		47: z5 <= -16'd100;
		48: z5 <= 16'd53;
		49: z5 <= 16'd71;
		50: z5 <= -16'd63;
		51: z5 <= 16'd102;
		52: z5 <= 16'd67;
		53: z5 <= 16'd124;
		54: z5 <= 16'd58;
		55: z5 <= -16'd89;
		56: z5 <= 16'd70;
		57: z5 <= -16'd3;
		58: z5 <= 16'd61;
		59: z5 <= 16'd89;
		60: z5 <= 16'd108;
		61: z5 <= -16'd97;
		62: z5 <= 16'd100;
		63: z5 <= -16'd62;
		64: z5 <= 16'd18;
		65: z5 <= 16'd96;
		66: z5 <= -16'd104;
		67: z5 <= 16'd0;
		68: z5 <= 16'd4;
		69: z5 <= -16'd110;
		70: z5 <= 16'd89;
		71: z5 <= -16'd20;
		72: z5 <= -16'd44;
		73: z5 <= 16'd78;
		74: z5 <= 16'd106;
		75: z5 <= 16'd96;
		76: z5 <= -16'd86;
		77: z5 <= -16'd76;
		78: z5 <= 16'd124;
		79: z5 <= 16'd96;
		80: z5 <= 16'd124;
		81: z5 <= -16'd67;
		82: z5 <= 16'd70;
		83: z5 <= 16'd63;
		84: z5 <= -16'd71;
		85: z5 <= 16'd0;
		86: z5 <= 16'd102;
		87: z5 <= 16'd127;
		88: z5 <= 16'd126;
		89: z5 <= 16'd35;
		90: z5 <= 16'd89;
		91: z5 <= 16'd106;
		92: z5 <= 16'd66;
		93: z5 <= 16'd61;
		94: z5 <= -16'd84;
		95: z5 <= -16'd43;
		96: z5 <= 16'd29;
		97: z5 <= -16'd60;
		98: z5 <= 16'd85;
		99: z5 <= -16'd94;
		100: z5 <= -16'd41;
		101: z5 <= 16'd46;
		102: z5 <= 16'd14;
		103: z5 <= 16'd43;
		104: z5 <= -16'd4;
		105: z5 <= -16'd8;
		106: z5 <= 16'd11;
		107: z5 <= 16'd39;
		108: z5 <= 16'd45;
		109: z5 <= 16'd8;
		110: z5 <= 16'd7;
		111: z5 <= 16'd41;
		112: z5 <= 16'd69;
		113: z5 <= -16'd51;
		114: z5 <= -16'd24;
		115: z5 <= 16'd127;
		116: z5 <= 16'd78;
		117: z5 <= -16'd50;
		118: z5 <= 16'd126;
		119: z5 <= 16'd76;
		120: z5 <= 16'd114;
		121: z5 <= 16'd87;
		122: z5 <= 16'd54;
		123: z5 <= 16'd52;
		124: z5 <= 16'd20;
		125: z5 <= 16'd98;
		126: z5 <= -16'd119;
		127: z5 <= -16'd78;
		endcase
		case(addr6)
		0: z6 <= 16'd119;
		1: z6 <= 16'd104;
		2: z6 <= -16'd111;
		3: z6 <= 16'd114;
		4: z6 <= -16'd1;
		5: z6 <= -16'd6;
		6: z6 <= 16'd39;
		7: z6 <= -16'd91;
		8: z6 <= -16'd21;
		9: z6 <= -16'd60;
		10: z6 <= -16'd57;
		11: z6 <= 16'd28;
		12: z6 <= 16'd21;
		13: z6 <= -16'd55;
		14: z6 <= -16'd26;
		15: z6 <= 16'd77;
		16: z6 <= 16'd17;
		17: z6 <= -16'd39;
		18: z6 <= -16'd3;
		19: z6 <= -16'd92;
		20: z6 <= -16'd79;
		21: z6 <= 16'd123;
		22: z6 <= 16'd59;
		23: z6 <= 16'd83;
		24: z6 <= -16'd28;
		25: z6 <= 16'd74;
		26: z6 <= 16'd67;
		27: z6 <= 16'd21;
		28: z6 <= -16'd109;
		29: z6 <= -16'd18;
		30: z6 <= -16'd30;
		31: z6 <= -16'd118;
		32: z6 <= -16'd42;
		33: z6 <= -16'd13;
		34: z6 <= 16'd124;
		35: z6 <= 16'd85;
		36: z6 <= 16'd109;
		37: z6 <= 16'd36;
		38: z6 <= 16'd122;
		39: z6 <= -16'd39;
		40: z6 <= 16'd104;
		41: z6 <= -16'd62;
		42: z6 <= 16'd117;
		43: z6 <= -16'd3;
		44: z6 <= 16'd11;
		45: z6 <= -16'd36;
		46: z6 <= -16'd54;
		47: z6 <= -16'd100;
		48: z6 <= 16'd53;
		49: z6 <= 16'd71;
		50: z6 <= -16'd63;
		51: z6 <= 16'd102;
		52: z6 <= 16'd67;
		53: z6 <= 16'd124;
		54: z6 <= 16'd58;
		55: z6 <= -16'd89;
		56: z6 <= 16'd70;
		57: z6 <= -16'd3;
		58: z6 <= 16'd61;
		59: z6 <= 16'd89;
		60: z6 <= 16'd108;
		61: z6 <= -16'd97;
		62: z6 <= 16'd100;
		63: z6 <= -16'd62;
		64: z6 <= 16'd18;
		65: z6 <= 16'd96;
		66: z6 <= -16'd104;
		67: z6 <= 16'd0;
		68: z6 <= 16'd4;
		69: z6 <= -16'd110;
		70: z6 <= 16'd89;
		71: z6 <= -16'd20;
		72: z6 <= -16'd44;
		73: z6 <= 16'd78;
		74: z6 <= 16'd106;
		75: z6 <= 16'd96;
		76: z6 <= -16'd86;
		77: z6 <= -16'd76;
		78: z6 <= 16'd124;
		79: z6 <= 16'd96;
		80: z6 <= 16'd124;
		81: z6 <= -16'd67;
		82: z6 <= 16'd70;
		83: z6 <= 16'd63;
		84: z6 <= -16'd71;
		85: z6 <= 16'd0;
		86: z6 <= 16'd102;
		87: z6 <= 16'd127;
		88: z6 <= 16'd126;
		89: z6 <= 16'd35;
		90: z6 <= 16'd89;
		91: z6 <= 16'd106;
		92: z6 <= 16'd66;
		93: z6 <= 16'd61;
		94: z6 <= -16'd84;
		95: z6 <= -16'd43;
		96: z6 <= 16'd29;
		97: z6 <= -16'd60;
		98: z6 <= 16'd85;
		99: z6 <= -16'd94;
		100: z6 <= -16'd41;
		101: z6 <= 16'd46;
		102: z6 <= 16'd14;
		103: z6 <= 16'd43;
		104: z6 <= -16'd4;
		105: z6 <= -16'd8;
		106: z6 <= 16'd11;
		107: z6 <= 16'd39;
		108: z6 <= 16'd45;
		109: z6 <= 16'd8;
		110: z6 <= 16'd7;
		111: z6 <= 16'd41;
		112: z6 <= 16'd69;
		113: z6 <= -16'd51;
		114: z6 <= -16'd24;
		115: z6 <= 16'd127;
		116: z6 <= 16'd78;
		117: z6 <= -16'd50;
		118: z6 <= 16'd126;
		119: z6 <= 16'd76;
		120: z6 <= 16'd114;
		121: z6 <= 16'd87;
		122: z6 <= 16'd54;
		123: z6 <= 16'd52;
		124: z6 <= 16'd20;
		125: z6 <= 16'd98;
		126: z6 <= -16'd119;
		127: z6 <= -16'd78;
		endcase
		case(addr7)
		0: z7 <= 16'd119;
		1: z7 <= 16'd104;
		2: z7 <= -16'd111;
		3: z7 <= 16'd114;
		4: z7 <= -16'd1;
		5: z7 <= -16'd6;
		6: z7 <= 16'd39;
		7: z7 <= -16'd91;
		8: z7 <= -16'd21;
		9: z7 <= -16'd60;
		10: z7 <= -16'd57;
		11: z7 <= 16'd28;
		12: z7 <= 16'd21;
		13: z7 <= -16'd55;
		14: z7 <= -16'd26;
		15: z7 <= 16'd77;
		16: z7 <= 16'd17;
		17: z7 <= -16'd39;
		18: z7 <= -16'd3;
		19: z7 <= -16'd92;
		20: z7 <= -16'd79;
		21: z7 <= 16'd123;
		22: z7 <= 16'd59;
		23: z7 <= 16'd83;
		24: z7 <= -16'd28;
		25: z7 <= 16'd74;
		26: z7 <= 16'd67;
		27: z7 <= 16'd21;
		28: z7 <= -16'd109;
		29: z7 <= -16'd18;
		30: z7 <= -16'd30;
		31: z7 <= -16'd118;
		32: z7 <= -16'd42;
		33: z7 <= -16'd13;
		34: z7 <= 16'd124;
		35: z7 <= 16'd85;
		36: z7 <= 16'd109;
		37: z7 <= 16'd36;
		38: z7 <= 16'd122;
		39: z7 <= -16'd39;
		40: z7 <= 16'd104;
		41: z7 <= -16'd62;
		42: z7 <= 16'd117;
		43: z7 <= -16'd3;
		44: z7 <= 16'd11;
		45: z7 <= -16'd36;
		46: z7 <= -16'd54;
		47: z7 <= -16'd100;
		48: z7 <= 16'd53;
		49: z7 <= 16'd71;
		50: z7 <= -16'd63;
		51: z7 <= 16'd102;
		52: z7 <= 16'd67;
		53: z7 <= 16'd124;
		54: z7 <= 16'd58;
		55: z7 <= -16'd89;
		56: z7 <= 16'd70;
		57: z7 <= -16'd3;
		58: z7 <= 16'd61;
		59: z7 <= 16'd89;
		60: z7 <= 16'd108;
		61: z7 <= -16'd97;
		62: z7 <= 16'd100;
		63: z7 <= -16'd62;
		64: z7 <= 16'd18;
		65: z7 <= 16'd96;
		66: z7 <= -16'd104;
		67: z7 <= 16'd0;
		68: z7 <= 16'd4;
		69: z7 <= -16'd110;
		70: z7 <= 16'd89;
		71: z7 <= -16'd20;
		72: z7 <= -16'd44;
		73: z7 <= 16'd78;
		74: z7 <= 16'd106;
		75: z7 <= 16'd96;
		76: z7 <= -16'd86;
		77: z7 <= -16'd76;
		78: z7 <= 16'd124;
		79: z7 <= 16'd96;
		80: z7 <= 16'd124;
		81: z7 <= -16'd67;
		82: z7 <= 16'd70;
		83: z7 <= 16'd63;
		84: z7 <= -16'd71;
		85: z7 <= 16'd0;
		86: z7 <= 16'd102;
		87: z7 <= 16'd127;
		88: z7 <= 16'd126;
		89: z7 <= 16'd35;
		90: z7 <= 16'd89;
		91: z7 <= 16'd106;
		92: z7 <= 16'd66;
		93: z7 <= 16'd61;
		94: z7 <= -16'd84;
		95: z7 <= -16'd43;
		96: z7 <= 16'd29;
		97: z7 <= -16'd60;
		98: z7 <= 16'd85;
		99: z7 <= -16'd94;
		100: z7 <= -16'd41;
		101: z7 <= 16'd46;
		102: z7 <= 16'd14;
		103: z7 <= 16'd43;
		104: z7 <= -16'd4;
		105: z7 <= -16'd8;
		106: z7 <= 16'd11;
		107: z7 <= 16'd39;
		108: z7 <= 16'd45;
		109: z7 <= 16'd8;
		110: z7 <= 16'd7;
		111: z7 <= 16'd41;
		112: z7 <= 16'd69;
		113: z7 <= -16'd51;
		114: z7 <= -16'd24;
		115: z7 <= 16'd127;
		116: z7 <= 16'd78;
		117: z7 <= -16'd50;
		118: z7 <= 16'd126;
		119: z7 <= 16'd76;
		120: z7 <= 16'd114;
		121: z7 <= 16'd87;
		122: z7 <= 16'd54;
		123: z7 <= 16'd52;
		124: z7 <= 16'd20;
		125: z7 <= 16'd98;
		126: z7 <= -16'd119;
		127: z7 <= -16'd78;
		endcase
	end
endmodule

