module fc_13_16_32_1_1(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 13;
	parameter N = 16;
	parameter T = 32;
	parameter R = 1;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned[7 : 0] addr_w;
	logic unsigned[3 : 0] addr_x;
	logic signed [31 : 0] v_out, m_out;
	logic unsigned wr_en_x;
	logic unsigned clear_acc;
	logic unsigned en_acc;

	controlFSM #(13,16) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr_w), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid));

	datapath #(32, 1) datapathMod(.clk(clk), .reset(reset), .m_out(m_out), .v_out(v_out),
									.en_acc(en_acc), .output_data(output_data), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	memory #(32, 16 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	fc_13_16_32_1_1_W_rom  matrixRom(.clk(clk), .addr(addr_w), .z(m_out));

endmodule

module fc_13_16_32_1_1_W_rom(clk, addr, z);
   input clk;
   input [7:0] addr;
   output logic signed [31:0] z;
   always_ff @(posedge clk) begin
      case(addr)
        0: z <= -32'd6370;
        1: z <= -32'd27204;
        2: z <= -32'd1490;
        3: z <= 32'd10299;
        4: z <= -32'd32735;
        5: z <= -32'd24362;
        6: z <= -32'd16502;
        7: z <= -32'd27717;
        8: z <= 32'd14015;
        9: z <= 32'd25893;
        10: z <= 32'd3385;
        11: z <= 32'd16193;
        12: z <= 32'd19209;
        13: z <= -32'd8654;
        14: z <= -32'd29767;
        15: z <= 32'd12507;
        16: z <= -32'd28465;
        17: z <= -32'd29370;
        18: z <= 32'd9207;
        19: z <= -32'd23541;
        20: z <= 32'd7627;
        21: z <= -32'd20947;
        22: z <= -32'd27771;
        23: z <= -32'd16077;
        24: z <= -32'd22555;
        25: z <= 32'd25622;
        26: z <= 32'd25772;
        27: z <= 32'd8993;
        28: z <= -32'd16559;
        29: z <= -32'd18548;
        30: z <= 32'd8074;
        31: z <= 32'd9839;
        32: z <= -32'd12983;
        33: z <= -32'd26184;
        34: z <= -32'd12630;
        35: z <= -32'd12950;
        36: z <= -32'd17778;
        37: z <= 32'd3636;
        38: z <= -32'd7899;
        39: z <= 32'd29006;
        40: z <= -32'd3239;
        41: z <= 32'd28254;
        42: z <= 32'd12431;
        43: z <= -32'd16798;
        44: z <= -32'd13168;
        45: z <= 32'd15432;
        46: z <= 32'd28477;
        47: z <= -32'd8865;
        48: z <= 32'd18831;
        49: z <= 32'd4916;
        50: z <= 32'd362;
        51: z <= -32'd6310;
        52: z <= 32'd16737;
        53: z <= 32'd5360;
        54: z <= 32'd10381;
        55: z <= 32'd26950;
        56: z <= -32'd1786;
        57: z <= 32'd3386;
        58: z <= 32'd3175;
        59: z <= 32'd14423;
        60: z <= 32'd17606;
        61: z <= -32'd21518;
        62: z <= -32'd8506;
        63: z <= -32'd28145;
        64: z <= -32'd14934;
        65: z <= 32'd11632;
        66: z <= -32'd8327;
        67: z <= 32'd57;
        68: z <= -32'd17500;
        69: z <= 32'd16542;
        70: z <= -32'd3705;
        71: z <= 32'd12030;
        72: z <= 32'd12029;
        73: z <= -32'd24042;
        74: z <= 32'd28000;
        75: z <= 32'd31629;
        76: z <= 32'd24159;
        77: z <= 32'd23710;
        78: z <= -32'd10003;
        79: z <= 32'd10222;
        80: z <= -32'd4142;
        81: z <= 32'd23127;
        82: z <= -32'd28856;
        83: z <= -32'd20172;
        84: z <= -32'd4281;
        85: z <= 32'd14294;
        86: z <= -32'd25990;
        87: z <= 32'd26701;
        88: z <= -32'd15088;
        89: z <= 32'd9954;
        90: z <= 32'd8356;
        91: z <= -32'd30250;
        92: z <= 32'd21204;
        93: z <= 32'd32618;
        94: z <= -32'd25626;
        95: z <= -32'd26498;
        96: z <= 32'd11482;
        97: z <= -32'd1185;
        98: z <= 32'd6327;
        99: z <= 32'd26751;
        100: z <= -32'd17410;
        101: z <= -32'd30146;
        102: z <= 32'd6013;
        103: z <= 32'd27387;
        104: z <= -32'd21419;
        105: z <= 32'd1245;
        106: z <= 32'd26248;
        107: z <= -32'd30028;
        108: z <= -32'd7813;
        109: z <= -32'd16523;
        110: z <= 32'd12962;
        111: z <= 32'd20814;
        112: z <= -32'd26163;
        113: z <= 32'd16874;
        114: z <= -32'd32126;
        115: z <= 32'd2324;
        116: z <= -32'd1600;
        117: z <= -32'd25348;
        118: z <= -32'd3742;
        119: z <= 32'd16080;
        120: z <= 32'd17374;
        121: z <= -32'd28154;
        122: z <= 32'd18599;
        123: z <= 32'd5810;
        124: z <= -32'd28303;
        125: z <= 32'd25741;
        126: z <= 32'd12081;
        127: z <= 32'd15947;
        128: z <= -32'd8212;
        129: z <= -32'd14360;
        130: z <= 32'd9930;
        131: z <= 32'd7146;
        132: z <= -32'd11737;
        133: z <= -32'd16825;
        134: z <= 32'd1765;
        135: z <= -32'd388;
        136: z <= 32'd17189;
        137: z <= -32'd4754;
        138: z <= 32'd2352;
        139: z <= -32'd23392;
        140: z <= 32'd11491;
        141: z <= -32'd17454;
        142: z <= 32'd30190;
        143: z <= 32'd18096;
        144: z <= 32'd32188;
        145: z <= 32'd30832;
        146: z <= -32'd12347;
        147: z <= -32'd2179;
        148: z <= -32'd27283;
        149: z <= 32'd16679;
        150: z <= -32'd18867;
        151: z <= 32'd22859;
        152: z <= 32'd21293;
        153: z <= 32'd32500;
        154: z <= -32'd4098;
        155: z <= 32'd25758;
        156: z <= 32'd25473;
        157: z <= -32'd24785;
        158: z <= 32'd8938;
        159: z <= -32'd15506;
        160: z <= -32'd6377;
        161: z <= -32'd13900;
        162: z <= 32'd24408;
        163: z <= 32'd14654;
        164: z <= 32'd2044;
        165: z <= -32'd6594;
        166: z <= -32'd18502;
        167: z <= -32'd13535;
        168: z <= 32'd21420;
        169: z <= 32'd16618;
        170: z <= -32'd4159;
        171: z <= 32'd143;
        172: z <= 32'd31932;
        173: z <= -32'd6736;
        174: z <= -32'd14528;
        175: z <= 32'd31353;
        176: z <= -32'd8672;
        177: z <= 32'd5893;
        178: z <= -32'd3594;
        179: z <= -32'd3187;
        180: z <= -32'd10196;
        181: z <= 32'd10307;
        182: z <= -32'd13095;
        183: z <= -32'd21671;
        184: z <= 32'd10040;
        185: z <= 32'd15575;
        186: z <= -32'd28680;
        187: z <= 32'd2745;
        188: z <= 32'd23558;
        189: z <= 32'd13026;
        190: z <= 32'd20007;
        191: z <= -32'd15587;
        192: z <= 32'd31894;
        193: z <= 32'd11648;
        194: z <= 32'd31836;
        195: z <= 32'd1170;
        196: z <= -32'd27714;
        197: z <= -32'd19434;
        198: z <= 32'd20403;
        199: z <= 32'd26474;
        200: z <= 32'd29953;
        201: z <= -32'd16523;
        202: z <= -32'd6151;
        203: z <= 32'd29117;
        204: z <= 32'd9509;
        205: z <= 32'd12089;
        206: z <= 32'd27702;
        207: z <= -32'd31931;
      endcase
   end
endmodule

