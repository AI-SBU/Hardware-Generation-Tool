`include "controlFSM.sv"
`include "datapath.sv"
`include "memory.sv"

module fc_16_8_16_1_4(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 16;
	parameter N = 8;
	parameter T = 16;
	parameter R = 1;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned [1 : 0] sel;

	logic signed [T-1 : 0] parallel_out0;
	logic signed [T-1 : 0] parallel_out1;
	logic signed [T-1 : 0] parallel_out2;
	logic signed [T-1 : 0] parallel_out3;

	logic unsigned[2 : 0] addr_x;
	logic signed [15 : 0] v_out;
	logic unsigned wr_en_x;

	logic unsigned[6 : 0] addr;

	logic unsigned[6 : 0] addr_w0;
	logic signed [15 : 0] m_out0;

	logic unsigned[6 : 0] addr_w1;
	logic signed [15 : 0] m_out1;

	logic unsigned[6 : 0] addr_w2;
	logic signed [15 : 0] m_out2;

	logic unsigned[6 : 0] addr_w3;
	logic signed [15 : 0] m_out3;

	logic unsigned clear_acc;
	logic unsigned en_acc;

	always_comb begin
		addr_w0 = addr + 0;
		addr_w1 = addr + 8;
		addr_w2 = addr + 16;
		addr_w3 = addr + 24;
	end

	controlFSM #(16,8,4) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid), .countToP(sel));

	memory #(16, 8 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	mux #(16, 4) muxMod(.parallel_out0(parallel_out0), .parallel_out1(parallel_out1), .parallel_out2(parallel_out2), .parallel_out3(parallel_out3), .sel(sel), .f(output_data));

	datapath #(16, 1) datapathMod0(.clk(clk), .reset(reset), .m_out(m_out0), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out0), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod1(.clk(clk), .reset(reset), .m_out(m_out1), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out1), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod2(.clk(clk), .reset(reset), .m_out(m_out2), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out2), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod3(.clk(clk), .reset(reset), .m_out(m_out3), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out3), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	fc_16_8_16_1_4_W_rom  matrixRom(.clk(clk),.addr0(addr_w0), .addr1(addr_w1), .addr2(addr_w2), .addr3(addr_w3), .z0(m_out0), .z1(m_out1), .z2(m_out2), .z3(m_out3));

endmodule

module mux(parallel_out0, parallel_out1, parallel_out2, parallel_out3, sel, f);
	parameter T = 16;
	parameter P = 4;

	output signed [T-1 : 0] f;
	input logic unsigned [1 : 0] sel;
	input signed [T-1 : 0] parallel_out0;
	input signed [T-1 : 0] parallel_out1;
	input signed [T-1 : 0] parallel_out2;
	input signed [T-1 : 0] parallel_out3;
	logic unsigned [P*T-1 : 0] array;
	assign  array = {parallel_out0[15 : 0], parallel_out1[15 : 0], parallel_out2[15 : 0], parallel_out3[15: 0]};

	assign f = (sel == 0) ? parallel_out0 : 
			(sel == 1) ? parallel_out1 : 
			(sel == 2) ? parallel_out2 : 
			(sel == 3) ? parallel_out3 : 16'bz;
endmodule

module fc_16_8_16_1_4_W_rom(clk, addr0, addr1, addr2, addr3, z0, z1, z2, z3);
	input clk;
	input [6:0] addr0;
	input [6:0] addr1;
	input [6:0] addr2;
	input [6:0] addr3;
	output logic signed [15:0] z0;
	output logic signed [15:0] z1;
	output logic signed [15:0] z2;
	output logic signed [15:0] z3;
	always_ff @(posedge clk) begin
		case(addr0)
		0: z0 <= -16'd115;
		1: z0 <= 16'd41;
		2: z0 <= -16'd73;
		3: z0 <= 16'd122;
		4: z0 <= 16'd110;
		5: z0 <= -16'd57;
		6: z0 <= -16'd119;
		7: z0 <= 16'd118;
		8: z0 <= -16'd111;
		9: z0 <= -16'd104;
		10: z0 <= -16'd52;
		11: z0 <= 16'd82;
		12: z0 <= -16'd103;
		13: z0 <= -16'd80;
		14: z0 <= -16'd91;
		15: z0 <= 16'd112;
		16: z0 <= 16'd18;
		17: z0 <= -16'd100;
		18: z0 <= 16'd79;
		19: z0 <= -16'd15;
		20: z0 <= -16'd58;
		21: z0 <= -16'd6;
		22: z0 <= -16'd124;
		23: z0 <= -16'd36;
		24: z0 <= -16'd83;
		25: z0 <= -16'd31;
		26: z0 <= -16'd97;
		27: z0 <= -16'd61;
		28: z0 <= -16'd39;
		29: z0 <= -16'd27;
		30: z0 <= 16'd119;
		31: z0 <= -16'd26;
		32: z0 <= -16'd114;
		33: z0 <= -16'd82;
		34: z0 <= -16'd32;
		35: z0 <= 16'd124;
		36: z0 <= -16'd10;
		37: z0 <= -16'd23;
		38: z0 <= 16'd114;
		39: z0 <= 16'd7;
		40: z0 <= 16'd1;
		41: z0 <= -16'd65;
		42: z0 <= -16'd38;
		43: z0 <= 16'd26;
		44: z0 <= -16'd17;
		45: z0 <= -16'd1;
		46: z0 <= 16'd11;
		47: z0 <= -16'd127;
		48: z0 <= 16'd28;
		49: z0 <= -16'd38;
		50: z0 <= -16'd14;
		51: z0 <= 16'd98;
		52: z0 <= 16'd85;
		53: z0 <= -16'd9;
		54: z0 <= -16'd66;
		55: z0 <= -16'd126;
		56: z0 <= 16'd88;
		57: z0 <= -16'd34;
		58: z0 <= -16'd59;
		59: z0 <= -16'd79;
		60: z0 <= 16'd67;
		61: z0 <= -16'd68;
		62: z0 <= 16'd23;
		63: z0 <= 16'd81;
		64: z0 <= -16'd21;
		65: z0 <= 16'd120;
		66: z0 <= 16'd77;
		67: z0 <= 16'd97;
		68: z0 <= -16'd31;
		69: z0 <= 16'd64;
		70: z0 <= -16'd24;
		71: z0 <= 16'd99;
		72: z0 <= 16'd127;
		73: z0 <= 16'd66;
		74: z0 <= -16'd3;
		75: z0 <= -16'd18;
		76: z0 <= -16'd62;
		77: z0 <= -16'd120;
		78: z0 <= -16'd17;
		79: z0 <= 16'd94;
		80: z0 <= -16'd29;
		81: z0 <= 16'd98;
		82: z0 <= 16'd64;
		83: z0 <= -16'd72;
		84: z0 <= -16'd39;
		85: z0 <= 16'd127;
		86: z0 <= -16'd70;
		87: z0 <= -16'd79;
		88: z0 <= -16'd35;
		89: z0 <= -16'd1;
		90: z0 <= -16'd29;
		91: z0 <= -16'd96;
		92: z0 <= 16'd59;
		93: z0 <= 16'd122;
		94: z0 <= 16'd113;
		95: z0 <= -16'd90;
		96: z0 <= 16'd114;
		97: z0 <= 16'd62;
		98: z0 <= -16'd121;
		99: z0 <= -16'd44;
		100: z0 <= -16'd2;
		101: z0 <= -16'd16;
		102: z0 <= -16'd73;
		103: z0 <= -16'd3;
		104: z0 <= -16'd78;
		105: z0 <= 16'd52;
		106: z0 <= 16'd107;
		107: z0 <= -16'd12;
		108: z0 <= 16'd61;
		109: z0 <= -16'd37;
		110: z0 <= -16'd46;
		111: z0 <= -16'd96;
		112: z0 <= -16'd67;
		113: z0 <= -16'd109;
		114: z0 <= -16'd40;
		115: z0 <= 16'd22;
		116: z0 <= -16'd110;
		117: z0 <= 16'd18;
		118: z0 <= 16'd71;
		119: z0 <= -16'd17;
		120: z0 <= -16'd111;
		121: z0 <= -16'd86;
		122: z0 <= 16'd15;
		123: z0 <= 16'd76;
		124: z0 <= -16'd91;
		125: z0 <= 16'd0;
		126: z0 <= 16'd115;
		127: z0 <= -16'd105;
		endcase
		case(addr1)
		0: z1 <= -16'd115;
		1: z1 <= 16'd41;
		2: z1 <= -16'd73;
		3: z1 <= 16'd122;
		4: z1 <= 16'd110;
		5: z1 <= -16'd57;
		6: z1 <= -16'd119;
		7: z1 <= 16'd118;
		8: z1 <= -16'd111;
		9: z1 <= -16'd104;
		10: z1 <= -16'd52;
		11: z1 <= 16'd82;
		12: z1 <= -16'd103;
		13: z1 <= -16'd80;
		14: z1 <= -16'd91;
		15: z1 <= 16'd112;
		16: z1 <= 16'd18;
		17: z1 <= -16'd100;
		18: z1 <= 16'd79;
		19: z1 <= -16'd15;
		20: z1 <= -16'd58;
		21: z1 <= -16'd6;
		22: z1 <= -16'd124;
		23: z1 <= -16'd36;
		24: z1 <= -16'd83;
		25: z1 <= -16'd31;
		26: z1 <= -16'd97;
		27: z1 <= -16'd61;
		28: z1 <= -16'd39;
		29: z1 <= -16'd27;
		30: z1 <= 16'd119;
		31: z1 <= -16'd26;
		32: z1 <= -16'd114;
		33: z1 <= -16'd82;
		34: z1 <= -16'd32;
		35: z1 <= 16'd124;
		36: z1 <= -16'd10;
		37: z1 <= -16'd23;
		38: z1 <= 16'd114;
		39: z1 <= 16'd7;
		40: z1 <= 16'd1;
		41: z1 <= -16'd65;
		42: z1 <= -16'd38;
		43: z1 <= 16'd26;
		44: z1 <= -16'd17;
		45: z1 <= -16'd1;
		46: z1 <= 16'd11;
		47: z1 <= -16'd127;
		48: z1 <= 16'd28;
		49: z1 <= -16'd38;
		50: z1 <= -16'd14;
		51: z1 <= 16'd98;
		52: z1 <= 16'd85;
		53: z1 <= -16'd9;
		54: z1 <= -16'd66;
		55: z1 <= -16'd126;
		56: z1 <= 16'd88;
		57: z1 <= -16'd34;
		58: z1 <= -16'd59;
		59: z1 <= -16'd79;
		60: z1 <= 16'd67;
		61: z1 <= -16'd68;
		62: z1 <= 16'd23;
		63: z1 <= 16'd81;
		64: z1 <= -16'd21;
		65: z1 <= 16'd120;
		66: z1 <= 16'd77;
		67: z1 <= 16'd97;
		68: z1 <= -16'd31;
		69: z1 <= 16'd64;
		70: z1 <= -16'd24;
		71: z1 <= 16'd99;
		72: z1 <= 16'd127;
		73: z1 <= 16'd66;
		74: z1 <= -16'd3;
		75: z1 <= -16'd18;
		76: z1 <= -16'd62;
		77: z1 <= -16'd120;
		78: z1 <= -16'd17;
		79: z1 <= 16'd94;
		80: z1 <= -16'd29;
		81: z1 <= 16'd98;
		82: z1 <= 16'd64;
		83: z1 <= -16'd72;
		84: z1 <= -16'd39;
		85: z1 <= 16'd127;
		86: z1 <= -16'd70;
		87: z1 <= -16'd79;
		88: z1 <= -16'd35;
		89: z1 <= -16'd1;
		90: z1 <= -16'd29;
		91: z1 <= -16'd96;
		92: z1 <= 16'd59;
		93: z1 <= 16'd122;
		94: z1 <= 16'd113;
		95: z1 <= -16'd90;
		96: z1 <= 16'd114;
		97: z1 <= 16'd62;
		98: z1 <= -16'd121;
		99: z1 <= -16'd44;
		100: z1 <= -16'd2;
		101: z1 <= -16'd16;
		102: z1 <= -16'd73;
		103: z1 <= -16'd3;
		104: z1 <= -16'd78;
		105: z1 <= 16'd52;
		106: z1 <= 16'd107;
		107: z1 <= -16'd12;
		108: z1 <= 16'd61;
		109: z1 <= -16'd37;
		110: z1 <= -16'd46;
		111: z1 <= -16'd96;
		112: z1 <= -16'd67;
		113: z1 <= -16'd109;
		114: z1 <= -16'd40;
		115: z1 <= 16'd22;
		116: z1 <= -16'd110;
		117: z1 <= 16'd18;
		118: z1 <= 16'd71;
		119: z1 <= -16'd17;
		120: z1 <= -16'd111;
		121: z1 <= -16'd86;
		122: z1 <= 16'd15;
		123: z1 <= 16'd76;
		124: z1 <= -16'd91;
		125: z1 <= 16'd0;
		126: z1 <= 16'd115;
		127: z1 <= -16'd105;
		endcase
		case(addr2)
		0: z2 <= -16'd115;
		1: z2 <= 16'd41;
		2: z2 <= -16'd73;
		3: z2 <= 16'd122;
		4: z2 <= 16'd110;
		5: z2 <= -16'd57;
		6: z2 <= -16'd119;
		7: z2 <= 16'd118;
		8: z2 <= -16'd111;
		9: z2 <= -16'd104;
		10: z2 <= -16'd52;
		11: z2 <= 16'd82;
		12: z2 <= -16'd103;
		13: z2 <= -16'd80;
		14: z2 <= -16'd91;
		15: z2 <= 16'd112;
		16: z2 <= 16'd18;
		17: z2 <= -16'd100;
		18: z2 <= 16'd79;
		19: z2 <= -16'd15;
		20: z2 <= -16'd58;
		21: z2 <= -16'd6;
		22: z2 <= -16'd124;
		23: z2 <= -16'd36;
		24: z2 <= -16'd83;
		25: z2 <= -16'd31;
		26: z2 <= -16'd97;
		27: z2 <= -16'd61;
		28: z2 <= -16'd39;
		29: z2 <= -16'd27;
		30: z2 <= 16'd119;
		31: z2 <= -16'd26;
		32: z2 <= -16'd114;
		33: z2 <= -16'd82;
		34: z2 <= -16'd32;
		35: z2 <= 16'd124;
		36: z2 <= -16'd10;
		37: z2 <= -16'd23;
		38: z2 <= 16'd114;
		39: z2 <= 16'd7;
		40: z2 <= 16'd1;
		41: z2 <= -16'd65;
		42: z2 <= -16'd38;
		43: z2 <= 16'd26;
		44: z2 <= -16'd17;
		45: z2 <= -16'd1;
		46: z2 <= 16'd11;
		47: z2 <= -16'd127;
		48: z2 <= 16'd28;
		49: z2 <= -16'd38;
		50: z2 <= -16'd14;
		51: z2 <= 16'd98;
		52: z2 <= 16'd85;
		53: z2 <= -16'd9;
		54: z2 <= -16'd66;
		55: z2 <= -16'd126;
		56: z2 <= 16'd88;
		57: z2 <= -16'd34;
		58: z2 <= -16'd59;
		59: z2 <= -16'd79;
		60: z2 <= 16'd67;
		61: z2 <= -16'd68;
		62: z2 <= 16'd23;
		63: z2 <= 16'd81;
		64: z2 <= -16'd21;
		65: z2 <= 16'd120;
		66: z2 <= 16'd77;
		67: z2 <= 16'd97;
		68: z2 <= -16'd31;
		69: z2 <= 16'd64;
		70: z2 <= -16'd24;
		71: z2 <= 16'd99;
		72: z2 <= 16'd127;
		73: z2 <= 16'd66;
		74: z2 <= -16'd3;
		75: z2 <= -16'd18;
		76: z2 <= -16'd62;
		77: z2 <= -16'd120;
		78: z2 <= -16'd17;
		79: z2 <= 16'd94;
		80: z2 <= -16'd29;
		81: z2 <= 16'd98;
		82: z2 <= 16'd64;
		83: z2 <= -16'd72;
		84: z2 <= -16'd39;
		85: z2 <= 16'd127;
		86: z2 <= -16'd70;
		87: z2 <= -16'd79;
		88: z2 <= -16'd35;
		89: z2 <= -16'd1;
		90: z2 <= -16'd29;
		91: z2 <= -16'd96;
		92: z2 <= 16'd59;
		93: z2 <= 16'd122;
		94: z2 <= 16'd113;
		95: z2 <= -16'd90;
		96: z2 <= 16'd114;
		97: z2 <= 16'd62;
		98: z2 <= -16'd121;
		99: z2 <= -16'd44;
		100: z2 <= -16'd2;
		101: z2 <= -16'd16;
		102: z2 <= -16'd73;
		103: z2 <= -16'd3;
		104: z2 <= -16'd78;
		105: z2 <= 16'd52;
		106: z2 <= 16'd107;
		107: z2 <= -16'd12;
		108: z2 <= 16'd61;
		109: z2 <= -16'd37;
		110: z2 <= -16'd46;
		111: z2 <= -16'd96;
		112: z2 <= -16'd67;
		113: z2 <= -16'd109;
		114: z2 <= -16'd40;
		115: z2 <= 16'd22;
		116: z2 <= -16'd110;
		117: z2 <= 16'd18;
		118: z2 <= 16'd71;
		119: z2 <= -16'd17;
		120: z2 <= -16'd111;
		121: z2 <= -16'd86;
		122: z2 <= 16'd15;
		123: z2 <= 16'd76;
		124: z2 <= -16'd91;
		125: z2 <= 16'd0;
		126: z2 <= 16'd115;
		127: z2 <= -16'd105;
		endcase
		case(addr3)
		0: z3 <= -16'd115;
		1: z3 <= 16'd41;
		2: z3 <= -16'd73;
		3: z3 <= 16'd122;
		4: z3 <= 16'd110;
		5: z3 <= -16'd57;
		6: z3 <= -16'd119;
		7: z3 <= 16'd118;
		8: z3 <= -16'd111;
		9: z3 <= -16'd104;
		10: z3 <= -16'd52;
		11: z3 <= 16'd82;
		12: z3 <= -16'd103;
		13: z3 <= -16'd80;
		14: z3 <= -16'd91;
		15: z3 <= 16'd112;
		16: z3 <= 16'd18;
		17: z3 <= -16'd100;
		18: z3 <= 16'd79;
		19: z3 <= -16'd15;
		20: z3 <= -16'd58;
		21: z3 <= -16'd6;
		22: z3 <= -16'd124;
		23: z3 <= -16'd36;
		24: z3 <= -16'd83;
		25: z3 <= -16'd31;
		26: z3 <= -16'd97;
		27: z3 <= -16'd61;
		28: z3 <= -16'd39;
		29: z3 <= -16'd27;
		30: z3 <= 16'd119;
		31: z3 <= -16'd26;
		32: z3 <= -16'd114;
		33: z3 <= -16'd82;
		34: z3 <= -16'd32;
		35: z3 <= 16'd124;
		36: z3 <= -16'd10;
		37: z3 <= -16'd23;
		38: z3 <= 16'd114;
		39: z3 <= 16'd7;
		40: z3 <= 16'd1;
		41: z3 <= -16'd65;
		42: z3 <= -16'd38;
		43: z3 <= 16'd26;
		44: z3 <= -16'd17;
		45: z3 <= -16'd1;
		46: z3 <= 16'd11;
		47: z3 <= -16'd127;
		48: z3 <= 16'd28;
		49: z3 <= -16'd38;
		50: z3 <= -16'd14;
		51: z3 <= 16'd98;
		52: z3 <= 16'd85;
		53: z3 <= -16'd9;
		54: z3 <= -16'd66;
		55: z3 <= -16'd126;
		56: z3 <= 16'd88;
		57: z3 <= -16'd34;
		58: z3 <= -16'd59;
		59: z3 <= -16'd79;
		60: z3 <= 16'd67;
		61: z3 <= -16'd68;
		62: z3 <= 16'd23;
		63: z3 <= 16'd81;
		64: z3 <= -16'd21;
		65: z3 <= 16'd120;
		66: z3 <= 16'd77;
		67: z3 <= 16'd97;
		68: z3 <= -16'd31;
		69: z3 <= 16'd64;
		70: z3 <= -16'd24;
		71: z3 <= 16'd99;
		72: z3 <= 16'd127;
		73: z3 <= 16'd66;
		74: z3 <= -16'd3;
		75: z3 <= -16'd18;
		76: z3 <= -16'd62;
		77: z3 <= -16'd120;
		78: z3 <= -16'd17;
		79: z3 <= 16'd94;
		80: z3 <= -16'd29;
		81: z3 <= 16'd98;
		82: z3 <= 16'd64;
		83: z3 <= -16'd72;
		84: z3 <= -16'd39;
		85: z3 <= 16'd127;
		86: z3 <= -16'd70;
		87: z3 <= -16'd79;
		88: z3 <= -16'd35;
		89: z3 <= -16'd1;
		90: z3 <= -16'd29;
		91: z3 <= -16'd96;
		92: z3 <= 16'd59;
		93: z3 <= 16'd122;
		94: z3 <= 16'd113;
		95: z3 <= -16'd90;
		96: z3 <= 16'd114;
		97: z3 <= 16'd62;
		98: z3 <= -16'd121;
		99: z3 <= -16'd44;
		100: z3 <= -16'd2;
		101: z3 <= -16'd16;
		102: z3 <= -16'd73;
		103: z3 <= -16'd3;
		104: z3 <= -16'd78;
		105: z3 <= 16'd52;
		106: z3 <= 16'd107;
		107: z3 <= -16'd12;
		108: z3 <= 16'd61;
		109: z3 <= -16'd37;
		110: z3 <= -16'd46;
		111: z3 <= -16'd96;
		112: z3 <= -16'd67;
		113: z3 <= -16'd109;
		114: z3 <= -16'd40;
		115: z3 <= 16'd22;
		116: z3 <= -16'd110;
		117: z3 <= 16'd18;
		118: z3 <= 16'd71;
		119: z3 <= -16'd17;
		120: z3 <= -16'd111;
		121: z3 <= -16'd86;
		122: z3 <= 16'd15;
		123: z3 <= 16'd76;
		124: z3 <= -16'd91;
		125: z3 <= 16'd0;
		126: z3 <= 16'd115;
		127: z3 <= -16'd105;
		endcase
	end
endmodule

