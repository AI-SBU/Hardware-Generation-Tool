`include "controlFSM.sv"
`include "datapath.sv"
`include "memory.sv"

module net_4_8_12_16_16_1_20(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);
	input clk, reset, input_valid, output_ready;
	input signed [15 : 0] input_data;
	output signed [15 : 0] output_data;
	output output_valid, input_ready;

	logic signed [15 : 0] layer1_output_data;
	logic unsigned layer1_output_valid;
	logic unsigned layer2_input_ready;
	logic signed [15 : 0] layer2_output_data;
	logic unsigned layer2_output_valid;
	logic unsigned layer3_input_ready;
   // this module should instantiate three layers and wire them together
l1_fc_8_4_16_1_4	layer1(.clk(clk), .reset(reset), .input_valid(input_valid), 
					.input_data(input_data), .input_ready(input_ready), .output_data(layer1_output_data), 
					.output_valid(layer1_output_valid), .output_ready(layer2_input_ready));
l2_fc_12_8_16_1_6	layer2(.clk(clk), .reset(reset), .input_data(layer1_output_data), .input_valid(layer1_output_valid), 
					 .input_ready(layer2_input_ready), .output_data(layer2_output_data), .output_valid(layer2_output_valid), .output_ready(layer3_input_ready));
l3_fc3_16_12_16_1_8	layer3(.clk(clk), .reset(reset), .input_data(layer2_output_data), .input_valid(layer2_output_valid), 
					 .input_ready(layer3_input_ready), .output_data(output_data), .output_valid(output_valid), .output_ready(output_ready));
endmodule

module l1_fc_8_4_16_1_4(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 8;
	parameter N = 4;
	parameter T = 16;
	parameter R = 1;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned [1 : 0] sel;

	logic signed [T-1 : 0] parallel_out0;
	logic signed [T-1 : 0] parallel_out1;
	logic signed [T-1 : 0] parallel_out2;
	logic signed [T-1 : 0] parallel_out3;

	logic unsigned[1 : 0] addr_x;
	logic signed [15 : 0] v_out;
	logic unsigned wr_en_x;

	logic unsigned[4 : 0] addr;

	logic unsigned[4 : 0] addr_w0;
	logic signed [15 : 0] m_out0;

	logic unsigned[4 : 0] addr_w1;
	logic signed [15 : 0] m_out1;

	logic unsigned[4 : 0] addr_w2;
	logic signed [15 : 0] m_out2;

	logic unsigned[4 : 0] addr_w3;
	logic signed [15 : 0] m_out3;

	logic unsigned clear_acc;
	logic unsigned en_acc;

	always_comb begin
		addr_w0 = addr + 0;
		addr_w1 = addr + 4;
		addr_w2 = addr + 8;
		addr_w3 = addr + 12;
	end

	controlFSM #(8,4,4) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid), .countToP(sel));

	memory #(16, 4 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	l1_fc_8_4_16_1_4_mux #(16, 4) muxMod(.parallel_out0(parallel_out0), .parallel_out1(parallel_out1), .parallel_out2(parallel_out2), .parallel_out3(parallel_out3), .sel(sel), .f(output_data));

	datapath #(16, 1) datapathMod0(.clk(clk), .reset(reset), .m_out(m_out0), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out0), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod1(.clk(clk), .reset(reset), .m_out(m_out1), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out1), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod2(.clk(clk), .reset(reset), .m_out(m_out2), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out2), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod3(.clk(clk), .reset(reset), .m_out(m_out3), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out3), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	l1_fc_8_4_16_1_4_W_rom  matrixRom(.clk(clk),.addr0(addr_w0), .addr1(addr_w1), .addr2(addr_w2), .addr3(addr_w3), .z0(m_out0), .z1(m_out1), .z2(m_out2), .z3(m_out3));

endmodule

module l1_fc_8_4_16_1_4_mux(parallel_out0, parallel_out1, parallel_out2, parallel_out3, sel, f);
	parameter T = 16;
	parameter P = 4;

	output signed [T-1 : 0] f;
	input logic unsigned [1 : 0] sel;
	input signed [T-1 : 0] parallel_out0;
	input signed [T-1 : 0] parallel_out1;
	input signed [T-1 : 0] parallel_out2;
	input signed [T-1 : 0] parallel_out3;
	logic unsigned [P*T-1 : 0] array;
	assign  array = {parallel_out0[15 : 0], parallel_out1[15 : 0], parallel_out2[15 : 0], parallel_out3[15: 0]};

	assign f = (sel == 0) ? parallel_out0 : 
			(sel == 1) ? parallel_out1 : 
			(sel == 2) ? parallel_out2 : 
			(sel == 3) ? parallel_out3 : 16'b0;
endmodule

module l1_fc_8_4_16_1_4_W_rom(clk, addr0, addr1, addr2, addr3, z0, z1, z2, z3);
	input clk;
	input [4:0] addr0;
	input [4:0] addr1;
	input [4:0] addr2;
	input [4:0] addr3;
	output logic signed [15:0] z0;
	output logic signed [15:0] z1;
	output logic signed [15:0] z2;
	output logic signed [15:0] z3;
	always_ff @(posedge clk) begin
		case(addr0)
		0: z0 <= 16'd5;
		1: z0 <= -16'd7;
		2: z0 <= 16'd0;
		3: z0 <= -16'd5;
		4: z0 <= -16'd5;
		5: z0 <= -16'd2;
		6: z0 <= -16'd7;
		7: z0 <= -16'd4;
		8: z0 <= 16'd3;
		9: z0 <= -16'd4;
		10: z0 <= -16'd1;
		11: z0 <= 16'd1;
		12: z0 <= 16'd5;
		13: z0 <= 16'd0;
		14: z0 <= 16'd2;
		15: z0 <= -16'd2;
		16: z0 <= 16'd5;
		17: z0 <= 16'd4;
		18: z0 <= 16'd2;
		19: z0 <= 16'd3;
		20: z0 <= 16'd7;
		21: z0 <= -16'd5;
		22: z0 <= -16'd1;
		23: z0 <= 16'd2;
		24: z0 <= -16'd7;
		25: z0 <= -16'd5;
		26: z0 <= -16'd2;
		27: z0 <= 16'd2;
		28: z0 <= -16'd5;
		29: z0 <= -16'd4;
		30: z0 <= -16'd3;
		31: z0 <= -16'd8;
		endcase
		case(addr1)
		0: z1 <= 16'd5;
		1: z1 <= -16'd7;
		2: z1 <= 16'd0;
		3: z1 <= -16'd5;
		4: z1 <= -16'd5;
		5: z1 <= -16'd2;
		6: z1 <= -16'd7;
		7: z1 <= -16'd4;
		8: z1 <= 16'd3;
		9: z1 <= -16'd4;
		10: z1 <= -16'd1;
		11: z1 <= 16'd1;
		12: z1 <= 16'd5;
		13: z1 <= 16'd0;
		14: z1 <= 16'd2;
		15: z1 <= -16'd2;
		16: z1 <= 16'd5;
		17: z1 <= 16'd4;
		18: z1 <= 16'd2;
		19: z1 <= 16'd3;
		20: z1 <= 16'd7;
		21: z1 <= -16'd5;
		22: z1 <= -16'd1;
		23: z1 <= 16'd2;
		24: z1 <= -16'd7;
		25: z1 <= -16'd5;
		26: z1 <= -16'd2;
		27: z1 <= 16'd2;
		28: z1 <= -16'd5;
		29: z1 <= -16'd4;
		30: z1 <= -16'd3;
		31: z1 <= -16'd8;
		endcase
		case(addr2)
		0: z2 <= 16'd5;
		1: z2 <= -16'd7;
		2: z2 <= 16'd0;
		3: z2 <= -16'd5;
		4: z2 <= -16'd5;
		5: z2 <= -16'd2;
		6: z2 <= -16'd7;
		7: z2 <= -16'd4;
		8: z2 <= 16'd3;
		9: z2 <= -16'd4;
		10: z2 <= -16'd1;
		11: z2 <= 16'd1;
		12: z2 <= 16'd5;
		13: z2 <= 16'd0;
		14: z2 <= 16'd2;
		15: z2 <= -16'd2;
		16: z2 <= 16'd5;
		17: z2 <= 16'd4;
		18: z2 <= 16'd2;
		19: z2 <= 16'd3;
		20: z2 <= 16'd7;
		21: z2 <= -16'd5;
		22: z2 <= -16'd1;
		23: z2 <= 16'd2;
		24: z2 <= -16'd7;
		25: z2 <= -16'd5;
		26: z2 <= -16'd2;
		27: z2 <= 16'd2;
		28: z2 <= -16'd5;
		29: z2 <= -16'd4;
		30: z2 <= -16'd3;
		31: z2 <= -16'd8;
		endcase
		case(addr3)
		0: z3 <= 16'd5;
		1: z3 <= -16'd7;
		2: z3 <= 16'd0;
		3: z3 <= -16'd5;
		4: z3 <= -16'd5;
		5: z3 <= -16'd2;
		6: z3 <= -16'd7;
		7: z3 <= -16'd4;
		8: z3 <= 16'd3;
		9: z3 <= -16'd4;
		10: z3 <= -16'd1;
		11: z3 <= 16'd1;
		12: z3 <= 16'd5;
		13: z3 <= 16'd0;
		14: z3 <= 16'd2;
		15: z3 <= -16'd2;
		16: z3 <= 16'd5;
		17: z3 <= 16'd4;
		18: z3 <= 16'd2;
		19: z3 <= 16'd3;
		20: z3 <= 16'd7;
		21: z3 <= -16'd5;
		22: z3 <= -16'd1;
		23: z3 <= 16'd2;
		24: z3 <= -16'd7;
		25: z3 <= -16'd5;
		26: z3 <= -16'd2;
		27: z3 <= 16'd2;
		28: z3 <= -16'd5;
		29: z3 <= -16'd4;
		30: z3 <= -16'd3;
		31: z3 <= -16'd8;
		endcase
	end
endmodule

module l2_fc_12_8_16_1_6(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 12;
	parameter N = 8;
	parameter T = 16;
	parameter R = 1;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned [2 : 0] sel;

	logic signed [T-1 : 0] parallel_out0;
	logic signed [T-1 : 0] parallel_out1;
	logic signed [T-1 : 0] parallel_out2;
	logic signed [T-1 : 0] parallel_out3;
	logic signed [T-1 : 0] parallel_out4;
	logic signed [T-1 : 0] parallel_out5;

	logic unsigned[2 : 0] addr_x;
	logic signed [15 : 0] v_out;
	logic unsigned wr_en_x;

	logic unsigned[6 : 0] addr;

	logic unsigned[6 : 0] addr_w0;
	logic signed [15 : 0] m_out0;

	logic unsigned[6 : 0] addr_w1;
	logic signed [15 : 0] m_out1;

	logic unsigned[6 : 0] addr_w2;
	logic signed [15 : 0] m_out2;

	logic unsigned[6 : 0] addr_w3;
	logic signed [15 : 0] m_out3;

	logic unsigned[6 : 0] addr_w4;
	logic signed [15 : 0] m_out4;

	logic unsigned[6 : 0] addr_w5;
	logic signed [15 : 0] m_out5;

	logic unsigned clear_acc;
	logic unsigned en_acc;

	always_comb begin
		addr_w0 = addr + 0;
		addr_w1 = addr + 8;
		addr_w2 = addr + 16;
		addr_w3 = addr + 24;
		addr_w4 = addr + 32;
		addr_w5 = addr + 40;
	end

	controlFSM #(12,8,6) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid), .countToP(sel));

	memory #(16, 8 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	l2_fc_12_8_16_1_6_mux #(16, 6) muxMod(.parallel_out0(parallel_out0), .parallel_out1(parallel_out1), .parallel_out2(parallel_out2), .parallel_out3(parallel_out3), .parallel_out4(parallel_out4), .parallel_out5(parallel_out5), .sel(sel), .f(output_data));

	datapath #(16, 1) datapathMod0(.clk(clk), .reset(reset), .m_out(m_out0), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out0), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod1(.clk(clk), .reset(reset), .m_out(m_out1), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out1), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod2(.clk(clk), .reset(reset), .m_out(m_out2), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out2), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod3(.clk(clk), .reset(reset), .m_out(m_out3), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out3), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod4(.clk(clk), .reset(reset), .m_out(m_out4), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out4), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod5(.clk(clk), .reset(reset), .m_out(m_out5), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out5), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	l2_fc_12_8_16_1_6_W_rom  matrixRom(.clk(clk),.addr0(addr_w0), .addr1(addr_w1), .addr2(addr_w2), .addr3(addr_w3), .addr4(addr_w4), .addr5(addr_w5), .z0(m_out0), .z1(m_out1), .z2(m_out2), .z3(m_out3), .z4(m_out4), .z5(m_out5));

endmodule

module l2_fc_12_8_16_1_6_mux(parallel_out0, parallel_out1, parallel_out2, parallel_out3, parallel_out4, parallel_out5, sel, f);
	parameter T = 16;
	parameter P = 6;

	output signed [T-1 : 0] f;
	input logic unsigned [2 : 0] sel;
	input signed [T-1 : 0] parallel_out0;
	input signed [T-1 : 0] parallel_out1;
	input signed [T-1 : 0] parallel_out2;
	input signed [T-1 : 0] parallel_out3;
	input signed [T-1 : 0] parallel_out4;
	input signed [T-1 : 0] parallel_out5;
	logic unsigned [P*T-1 : 0] array;
	assign  array = {parallel_out0[15 : 0], parallel_out1[15 : 0], parallel_out2[15 : 0], parallel_out3[15 : 0], parallel_out4[15 : 0], parallel_out5[15: 0]};

	assign f = (sel == 0) ? parallel_out0 : 
			(sel == 1) ? parallel_out1 : 
			(sel == 2) ? parallel_out2 : 
			(sel == 3) ? parallel_out3 : 
			(sel == 4) ? parallel_out4 : 
			(sel == 5) ? parallel_out5 : 16'b0;
endmodule

module l2_fc_12_8_16_1_6_W_rom(clk, addr0, addr1, addr2, addr3, addr4, addr5, z0, z1, z2, z3, z4, z5);
	input clk;
	input [6:0] addr0;
	input [6:0] addr1;
	input [6:0] addr2;
	input [6:0] addr3;
	input [6:0] addr4;
	input [6:0] addr5;
	output logic signed [15:0] z0;
	output logic signed [15:0] z1;
	output logic signed [15:0] z2;
	output logic signed [15:0] z3;
	output logic signed [15:0] z4;
	output logic signed [15:0] z5;
	always_ff @(posedge clk) begin
		case(addr0)
		0: z0 <= -16'd2;
		1: z0 <= 16'd5;
		2: z0 <= -16'd5;
		3: z0 <= 16'd1;
		4: z0 <= -16'd4;
		5: z0 <= -16'd4;
		6: z0 <= 16'd5;
		7: z0 <= 16'd7;
		8: z0 <= 16'd0;
		9: z0 <= -16'd4;
		10: z0 <= 16'd0;
		11: z0 <= -16'd2;
		12: z0 <= 16'd5;
		13: z0 <= -16'd6;
		14: z0 <= 16'd4;
		15: z0 <= 16'd2;
		16: z0 <= 16'd6;
		17: z0 <= -16'd2;
		18: z0 <= -16'd2;
		19: z0 <= 16'd6;
		20: z0 <= 16'd1;
		21: z0 <= 16'd5;
		22: z0 <= 16'd0;
		23: z0 <= 16'd3;
		24: z0 <= -16'd8;
		25: z0 <= 16'd6;
		26: z0 <= -16'd3;
		27: z0 <= -16'd5;
		28: z0 <= -16'd6;
		29: z0 <= 16'd2;
		30: z0 <= -16'd5;
		31: z0 <= 16'd0;
		32: z0 <= -16'd1;
		33: z0 <= -16'd2;
		34: z0 <= -16'd6;
		35: z0 <= 16'd3;
		36: z0 <= 16'd2;
		37: z0 <= 16'd7;
		38: z0 <= 16'd2;
		39: z0 <= -16'd6;
		40: z0 <= -16'd4;
		41: z0 <= -16'd5;
		42: z0 <= 16'd0;
		43: z0 <= -16'd7;
		44: z0 <= -16'd3;
		45: z0 <= -16'd4;
		46: z0 <= 16'd3;
		47: z0 <= -16'd4;
		48: z0 <= 16'd3;
		49: z0 <= -16'd7;
		50: z0 <= -16'd6;
		51: z0 <= -16'd4;
		52: z0 <= 16'd6;
		53: z0 <= 16'd2;
		54: z0 <= 16'd7;
		55: z0 <= 16'd6;
		56: z0 <= 16'd0;
		57: z0 <= -16'd4;
		58: z0 <= -16'd7;
		59: z0 <= 16'd2;
		60: z0 <= 16'd6;
		61: z0 <= -16'd4;
		62: z0 <= -16'd5;
		63: z0 <= -16'd2;
		64: z0 <= 16'd2;
		65: z0 <= -16'd3;
		66: z0 <= -16'd7;
		67: z0 <= -16'd4;
		68: z0 <= -16'd4;
		69: z0 <= 16'd4;
		70: z0 <= -16'd1;
		71: z0 <= 16'd0;
		72: z0 <= 16'd7;
		73: z0 <= 16'd7;
		74: z0 <= 16'd1;
		75: z0 <= -16'd4;
		76: z0 <= -16'd4;
		77: z0 <= -16'd3;
		78: z0 <= 16'd0;
		79: z0 <= 16'd7;
		80: z0 <= -16'd2;
		81: z0 <= 16'd2;
		82: z0 <= -16'd5;
		83: z0 <= -16'd3;
		84: z0 <= -16'd4;
		85: z0 <= -16'd5;
		86: z0 <= -16'd5;
		87: z0 <= 16'd4;
		88: z0 <= -16'd1;
		89: z0 <= -16'd3;
		90: z0 <= -16'd1;
		91: z0 <= -16'd2;
		92: z0 <= 16'd1;
		93: z0 <= 16'd2;
		94: z0 <= 16'd4;
		95: z0 <= -16'd4;
		endcase
		case(addr1)
		0: z1 <= -16'd2;
		1: z1 <= 16'd5;
		2: z1 <= -16'd5;
		3: z1 <= 16'd1;
		4: z1 <= -16'd4;
		5: z1 <= -16'd4;
		6: z1 <= 16'd5;
		7: z1 <= 16'd7;
		8: z1 <= 16'd0;
		9: z1 <= -16'd4;
		10: z1 <= 16'd0;
		11: z1 <= -16'd2;
		12: z1 <= 16'd5;
		13: z1 <= -16'd6;
		14: z1 <= 16'd4;
		15: z1 <= 16'd2;
		16: z1 <= 16'd6;
		17: z1 <= -16'd2;
		18: z1 <= -16'd2;
		19: z1 <= 16'd6;
		20: z1 <= 16'd1;
		21: z1 <= 16'd5;
		22: z1 <= 16'd0;
		23: z1 <= 16'd3;
		24: z1 <= -16'd8;
		25: z1 <= 16'd6;
		26: z1 <= -16'd3;
		27: z1 <= -16'd5;
		28: z1 <= -16'd6;
		29: z1 <= 16'd2;
		30: z1 <= -16'd5;
		31: z1 <= 16'd0;
		32: z1 <= -16'd1;
		33: z1 <= -16'd2;
		34: z1 <= -16'd6;
		35: z1 <= 16'd3;
		36: z1 <= 16'd2;
		37: z1 <= 16'd7;
		38: z1 <= 16'd2;
		39: z1 <= -16'd6;
		40: z1 <= -16'd4;
		41: z1 <= -16'd5;
		42: z1 <= 16'd0;
		43: z1 <= -16'd7;
		44: z1 <= -16'd3;
		45: z1 <= -16'd4;
		46: z1 <= 16'd3;
		47: z1 <= -16'd4;
		48: z1 <= 16'd3;
		49: z1 <= -16'd7;
		50: z1 <= -16'd6;
		51: z1 <= -16'd4;
		52: z1 <= 16'd6;
		53: z1 <= 16'd2;
		54: z1 <= 16'd7;
		55: z1 <= 16'd6;
		56: z1 <= 16'd0;
		57: z1 <= -16'd4;
		58: z1 <= -16'd7;
		59: z1 <= 16'd2;
		60: z1 <= 16'd6;
		61: z1 <= -16'd4;
		62: z1 <= -16'd5;
		63: z1 <= -16'd2;
		64: z1 <= 16'd2;
		65: z1 <= -16'd3;
		66: z1 <= -16'd7;
		67: z1 <= -16'd4;
		68: z1 <= -16'd4;
		69: z1 <= 16'd4;
		70: z1 <= -16'd1;
		71: z1 <= 16'd0;
		72: z1 <= 16'd7;
		73: z1 <= 16'd7;
		74: z1 <= 16'd1;
		75: z1 <= -16'd4;
		76: z1 <= -16'd4;
		77: z1 <= -16'd3;
		78: z1 <= 16'd0;
		79: z1 <= 16'd7;
		80: z1 <= -16'd2;
		81: z1 <= 16'd2;
		82: z1 <= -16'd5;
		83: z1 <= -16'd3;
		84: z1 <= -16'd4;
		85: z1 <= -16'd5;
		86: z1 <= -16'd5;
		87: z1 <= 16'd4;
		88: z1 <= -16'd1;
		89: z1 <= -16'd3;
		90: z1 <= -16'd1;
		91: z1 <= -16'd2;
		92: z1 <= 16'd1;
		93: z1 <= 16'd2;
		94: z1 <= 16'd4;
		95: z1 <= -16'd4;
		endcase
		case(addr2)
		0: z2 <= -16'd2;
		1: z2 <= 16'd5;
		2: z2 <= -16'd5;
		3: z2 <= 16'd1;
		4: z2 <= -16'd4;
		5: z2 <= -16'd4;
		6: z2 <= 16'd5;
		7: z2 <= 16'd7;
		8: z2 <= 16'd0;
		9: z2 <= -16'd4;
		10: z2 <= 16'd0;
		11: z2 <= -16'd2;
		12: z2 <= 16'd5;
		13: z2 <= -16'd6;
		14: z2 <= 16'd4;
		15: z2 <= 16'd2;
		16: z2 <= 16'd6;
		17: z2 <= -16'd2;
		18: z2 <= -16'd2;
		19: z2 <= 16'd6;
		20: z2 <= 16'd1;
		21: z2 <= 16'd5;
		22: z2 <= 16'd0;
		23: z2 <= 16'd3;
		24: z2 <= -16'd8;
		25: z2 <= 16'd6;
		26: z2 <= -16'd3;
		27: z2 <= -16'd5;
		28: z2 <= -16'd6;
		29: z2 <= 16'd2;
		30: z2 <= -16'd5;
		31: z2 <= 16'd0;
		32: z2 <= -16'd1;
		33: z2 <= -16'd2;
		34: z2 <= -16'd6;
		35: z2 <= 16'd3;
		36: z2 <= 16'd2;
		37: z2 <= 16'd7;
		38: z2 <= 16'd2;
		39: z2 <= -16'd6;
		40: z2 <= -16'd4;
		41: z2 <= -16'd5;
		42: z2 <= 16'd0;
		43: z2 <= -16'd7;
		44: z2 <= -16'd3;
		45: z2 <= -16'd4;
		46: z2 <= 16'd3;
		47: z2 <= -16'd4;
		48: z2 <= 16'd3;
		49: z2 <= -16'd7;
		50: z2 <= -16'd6;
		51: z2 <= -16'd4;
		52: z2 <= 16'd6;
		53: z2 <= 16'd2;
		54: z2 <= 16'd7;
		55: z2 <= 16'd6;
		56: z2 <= 16'd0;
		57: z2 <= -16'd4;
		58: z2 <= -16'd7;
		59: z2 <= 16'd2;
		60: z2 <= 16'd6;
		61: z2 <= -16'd4;
		62: z2 <= -16'd5;
		63: z2 <= -16'd2;
		64: z2 <= 16'd2;
		65: z2 <= -16'd3;
		66: z2 <= -16'd7;
		67: z2 <= -16'd4;
		68: z2 <= -16'd4;
		69: z2 <= 16'd4;
		70: z2 <= -16'd1;
		71: z2 <= 16'd0;
		72: z2 <= 16'd7;
		73: z2 <= 16'd7;
		74: z2 <= 16'd1;
		75: z2 <= -16'd4;
		76: z2 <= -16'd4;
		77: z2 <= -16'd3;
		78: z2 <= 16'd0;
		79: z2 <= 16'd7;
		80: z2 <= -16'd2;
		81: z2 <= 16'd2;
		82: z2 <= -16'd5;
		83: z2 <= -16'd3;
		84: z2 <= -16'd4;
		85: z2 <= -16'd5;
		86: z2 <= -16'd5;
		87: z2 <= 16'd4;
		88: z2 <= -16'd1;
		89: z2 <= -16'd3;
		90: z2 <= -16'd1;
		91: z2 <= -16'd2;
		92: z2 <= 16'd1;
		93: z2 <= 16'd2;
		94: z2 <= 16'd4;
		95: z2 <= -16'd4;
		endcase
		case(addr3)
		0: z3 <= -16'd2;
		1: z3 <= 16'd5;
		2: z3 <= -16'd5;
		3: z3 <= 16'd1;
		4: z3 <= -16'd4;
		5: z3 <= -16'd4;
		6: z3 <= 16'd5;
		7: z3 <= 16'd7;
		8: z3 <= 16'd0;
		9: z3 <= -16'd4;
		10: z3 <= 16'd0;
		11: z3 <= -16'd2;
		12: z3 <= 16'd5;
		13: z3 <= -16'd6;
		14: z3 <= 16'd4;
		15: z3 <= 16'd2;
		16: z3 <= 16'd6;
		17: z3 <= -16'd2;
		18: z3 <= -16'd2;
		19: z3 <= 16'd6;
		20: z3 <= 16'd1;
		21: z3 <= 16'd5;
		22: z3 <= 16'd0;
		23: z3 <= 16'd3;
		24: z3 <= -16'd8;
		25: z3 <= 16'd6;
		26: z3 <= -16'd3;
		27: z3 <= -16'd5;
		28: z3 <= -16'd6;
		29: z3 <= 16'd2;
		30: z3 <= -16'd5;
		31: z3 <= 16'd0;
		32: z3 <= -16'd1;
		33: z3 <= -16'd2;
		34: z3 <= -16'd6;
		35: z3 <= 16'd3;
		36: z3 <= 16'd2;
		37: z3 <= 16'd7;
		38: z3 <= 16'd2;
		39: z3 <= -16'd6;
		40: z3 <= -16'd4;
		41: z3 <= -16'd5;
		42: z3 <= 16'd0;
		43: z3 <= -16'd7;
		44: z3 <= -16'd3;
		45: z3 <= -16'd4;
		46: z3 <= 16'd3;
		47: z3 <= -16'd4;
		48: z3 <= 16'd3;
		49: z3 <= -16'd7;
		50: z3 <= -16'd6;
		51: z3 <= -16'd4;
		52: z3 <= 16'd6;
		53: z3 <= 16'd2;
		54: z3 <= 16'd7;
		55: z3 <= 16'd6;
		56: z3 <= 16'd0;
		57: z3 <= -16'd4;
		58: z3 <= -16'd7;
		59: z3 <= 16'd2;
		60: z3 <= 16'd6;
		61: z3 <= -16'd4;
		62: z3 <= -16'd5;
		63: z3 <= -16'd2;
		64: z3 <= 16'd2;
		65: z3 <= -16'd3;
		66: z3 <= -16'd7;
		67: z3 <= -16'd4;
		68: z3 <= -16'd4;
		69: z3 <= 16'd4;
		70: z3 <= -16'd1;
		71: z3 <= 16'd0;
		72: z3 <= 16'd7;
		73: z3 <= 16'd7;
		74: z3 <= 16'd1;
		75: z3 <= -16'd4;
		76: z3 <= -16'd4;
		77: z3 <= -16'd3;
		78: z3 <= 16'd0;
		79: z3 <= 16'd7;
		80: z3 <= -16'd2;
		81: z3 <= 16'd2;
		82: z3 <= -16'd5;
		83: z3 <= -16'd3;
		84: z3 <= -16'd4;
		85: z3 <= -16'd5;
		86: z3 <= -16'd5;
		87: z3 <= 16'd4;
		88: z3 <= -16'd1;
		89: z3 <= -16'd3;
		90: z3 <= -16'd1;
		91: z3 <= -16'd2;
		92: z3 <= 16'd1;
		93: z3 <= 16'd2;
		94: z3 <= 16'd4;
		95: z3 <= -16'd4;
		endcase
		case(addr4)
		0: z4 <= -16'd2;
		1: z4 <= 16'd5;
		2: z4 <= -16'd5;
		3: z4 <= 16'd1;
		4: z4 <= -16'd4;
		5: z4 <= -16'd4;
		6: z4 <= 16'd5;
		7: z4 <= 16'd7;
		8: z4 <= 16'd0;
		9: z4 <= -16'd4;
		10: z4 <= 16'd0;
		11: z4 <= -16'd2;
		12: z4 <= 16'd5;
		13: z4 <= -16'd6;
		14: z4 <= 16'd4;
		15: z4 <= 16'd2;
		16: z4 <= 16'd6;
		17: z4 <= -16'd2;
		18: z4 <= -16'd2;
		19: z4 <= 16'd6;
		20: z4 <= 16'd1;
		21: z4 <= 16'd5;
		22: z4 <= 16'd0;
		23: z4 <= 16'd3;
		24: z4 <= -16'd8;
		25: z4 <= 16'd6;
		26: z4 <= -16'd3;
		27: z4 <= -16'd5;
		28: z4 <= -16'd6;
		29: z4 <= 16'd2;
		30: z4 <= -16'd5;
		31: z4 <= 16'd0;
		32: z4 <= -16'd1;
		33: z4 <= -16'd2;
		34: z4 <= -16'd6;
		35: z4 <= 16'd3;
		36: z4 <= 16'd2;
		37: z4 <= 16'd7;
		38: z4 <= 16'd2;
		39: z4 <= -16'd6;
		40: z4 <= -16'd4;
		41: z4 <= -16'd5;
		42: z4 <= 16'd0;
		43: z4 <= -16'd7;
		44: z4 <= -16'd3;
		45: z4 <= -16'd4;
		46: z4 <= 16'd3;
		47: z4 <= -16'd4;
		48: z4 <= 16'd3;
		49: z4 <= -16'd7;
		50: z4 <= -16'd6;
		51: z4 <= -16'd4;
		52: z4 <= 16'd6;
		53: z4 <= 16'd2;
		54: z4 <= 16'd7;
		55: z4 <= 16'd6;
		56: z4 <= 16'd0;
		57: z4 <= -16'd4;
		58: z4 <= -16'd7;
		59: z4 <= 16'd2;
		60: z4 <= 16'd6;
		61: z4 <= -16'd4;
		62: z4 <= -16'd5;
		63: z4 <= -16'd2;
		64: z4 <= 16'd2;
		65: z4 <= -16'd3;
		66: z4 <= -16'd7;
		67: z4 <= -16'd4;
		68: z4 <= -16'd4;
		69: z4 <= 16'd4;
		70: z4 <= -16'd1;
		71: z4 <= 16'd0;
		72: z4 <= 16'd7;
		73: z4 <= 16'd7;
		74: z4 <= 16'd1;
		75: z4 <= -16'd4;
		76: z4 <= -16'd4;
		77: z4 <= -16'd3;
		78: z4 <= 16'd0;
		79: z4 <= 16'd7;
		80: z4 <= -16'd2;
		81: z4 <= 16'd2;
		82: z4 <= -16'd5;
		83: z4 <= -16'd3;
		84: z4 <= -16'd4;
		85: z4 <= -16'd5;
		86: z4 <= -16'd5;
		87: z4 <= 16'd4;
		88: z4 <= -16'd1;
		89: z4 <= -16'd3;
		90: z4 <= -16'd1;
		91: z4 <= -16'd2;
		92: z4 <= 16'd1;
		93: z4 <= 16'd2;
		94: z4 <= 16'd4;
		95: z4 <= -16'd4;
		endcase
		case(addr5)
		0: z5 <= -16'd2;
		1: z5 <= 16'd5;
		2: z5 <= -16'd5;
		3: z5 <= 16'd1;
		4: z5 <= -16'd4;
		5: z5 <= -16'd4;
		6: z5 <= 16'd5;
		7: z5 <= 16'd7;
		8: z5 <= 16'd0;
		9: z5 <= -16'd4;
		10: z5 <= 16'd0;
		11: z5 <= -16'd2;
		12: z5 <= 16'd5;
		13: z5 <= -16'd6;
		14: z5 <= 16'd4;
		15: z5 <= 16'd2;
		16: z5 <= 16'd6;
		17: z5 <= -16'd2;
		18: z5 <= -16'd2;
		19: z5 <= 16'd6;
		20: z5 <= 16'd1;
		21: z5 <= 16'd5;
		22: z5 <= 16'd0;
		23: z5 <= 16'd3;
		24: z5 <= -16'd8;
		25: z5 <= 16'd6;
		26: z5 <= -16'd3;
		27: z5 <= -16'd5;
		28: z5 <= -16'd6;
		29: z5 <= 16'd2;
		30: z5 <= -16'd5;
		31: z5 <= 16'd0;
		32: z5 <= -16'd1;
		33: z5 <= -16'd2;
		34: z5 <= -16'd6;
		35: z5 <= 16'd3;
		36: z5 <= 16'd2;
		37: z5 <= 16'd7;
		38: z5 <= 16'd2;
		39: z5 <= -16'd6;
		40: z5 <= -16'd4;
		41: z5 <= -16'd5;
		42: z5 <= 16'd0;
		43: z5 <= -16'd7;
		44: z5 <= -16'd3;
		45: z5 <= -16'd4;
		46: z5 <= 16'd3;
		47: z5 <= -16'd4;
		48: z5 <= 16'd3;
		49: z5 <= -16'd7;
		50: z5 <= -16'd6;
		51: z5 <= -16'd4;
		52: z5 <= 16'd6;
		53: z5 <= 16'd2;
		54: z5 <= 16'd7;
		55: z5 <= 16'd6;
		56: z5 <= 16'd0;
		57: z5 <= -16'd4;
		58: z5 <= -16'd7;
		59: z5 <= 16'd2;
		60: z5 <= 16'd6;
		61: z5 <= -16'd4;
		62: z5 <= -16'd5;
		63: z5 <= -16'd2;
		64: z5 <= 16'd2;
		65: z5 <= -16'd3;
		66: z5 <= -16'd7;
		67: z5 <= -16'd4;
		68: z5 <= -16'd4;
		69: z5 <= 16'd4;
		70: z5 <= -16'd1;
		71: z5 <= 16'd0;
		72: z5 <= 16'd7;
		73: z5 <= 16'd7;
		74: z5 <= 16'd1;
		75: z5 <= -16'd4;
		76: z5 <= -16'd4;
		77: z5 <= -16'd3;
		78: z5 <= 16'd0;
		79: z5 <= 16'd7;
		80: z5 <= -16'd2;
		81: z5 <= 16'd2;
		82: z5 <= -16'd5;
		83: z5 <= -16'd3;
		84: z5 <= -16'd4;
		85: z5 <= -16'd5;
		86: z5 <= -16'd5;
		87: z5 <= 16'd4;
		88: z5 <= -16'd1;
		89: z5 <= -16'd3;
		90: z5 <= -16'd1;
		91: z5 <= -16'd2;
		92: z5 <= 16'd1;
		93: z5 <= 16'd2;
		94: z5 <= 16'd4;
		95: z5 <= -16'd4;
		endcase
	end
endmodule

module l3_fc3_16_12_16_1_8(clk, reset, input_valid, input_ready, input_data, output_valid, output_ready, output_data);

	parameter M = 16;
	parameter N = 12;
	parameter T = 16;
	parameter R = 1;
	localparam LOGSIZE_M = $clog2(M*N);
	localparam LOGSIZE_N = $clog2(N);

	input clk, reset, input_valid, output_ready;
	input signed [T-1 : 0] input_data;
	output signed [T-1 : 0] output_data;
	output output_valid, input_ready;

	logic unsigned [2 : 0] sel;

	logic signed [T-1 : 0] parallel_out0;
	logic signed [T-1 : 0] parallel_out1;
	logic signed [T-1 : 0] parallel_out2;
	logic signed [T-1 : 0] parallel_out3;
	logic signed [T-1 : 0] parallel_out4;
	logic signed [T-1 : 0] parallel_out5;
	logic signed [T-1 : 0] parallel_out6;
	logic signed [T-1 : 0] parallel_out7;

	logic unsigned[3 : 0] addr_x;
	logic signed [15 : 0] v_out;
	logic unsigned wr_en_x;

	logic unsigned[7 : 0] addr;

	logic unsigned[7 : 0] addr_w0;
	logic signed [15 : 0] m_out0;

	logic unsigned[7 : 0] addr_w1;
	logic signed [15 : 0] m_out1;

	logic unsigned[7 : 0] addr_w2;
	logic signed [15 : 0] m_out2;

	logic unsigned[7 : 0] addr_w3;
	logic signed [15 : 0] m_out3;

	logic unsigned[7 : 0] addr_w4;
	logic signed [15 : 0] m_out4;

	logic unsigned[7 : 0] addr_w5;
	logic signed [15 : 0] m_out5;

	logic unsigned[7 : 0] addr_w6;
	logic signed [15 : 0] m_out6;

	logic unsigned[7 : 0] addr_w7;
	logic signed [15 : 0] m_out7;

	logic unsigned clear_acc;
	logic unsigned en_acc;

	always_comb begin
		addr_w0 = addr + 0;
		addr_w1 = addr + 12;
		addr_w2 = addr + 24;
		addr_w3 = addr + 36;
		addr_w4 = addr + 48;
		addr_w5 = addr + 60;
		addr_w6 = addr + 72;
		addr_w7 = addr + 84;
	end

	controlFSM #(16,12,8) controlMod(.clk(clk), .reset(reset), .input_valid(input_valid), .output_ready(output_ready),
									.addr_x(addr_x) , .wr_en_x(wr_en_x),.addr_w(addr), .en_acc(en_acc), .clear_acc(clear_acc),
									.input_ready(input_ready), .output_valid(output_valid), .countToP(sel));

	memory #(16, 12 )  vector(.clk(clk), .data_in(input_data), .data_out(v_out), .addr(addr_x), .wr_en(wr_en_x));

	l3_fc3_16_12_16_1_8_mux #(16, 8) muxMod(.parallel_out0(parallel_out0), .parallel_out1(parallel_out1), .parallel_out2(parallel_out2), .parallel_out3(parallel_out3), .parallel_out4(parallel_out4), .parallel_out5(parallel_out5), .parallel_out6(parallel_out6), .parallel_out7(parallel_out7), .sel(sel), .f(output_data));

	datapath #(16, 1) datapathMod0(.clk(clk), .reset(reset), .m_out(m_out0), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out0), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod1(.clk(clk), .reset(reset), .m_out(m_out1), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out1), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod2(.clk(clk), .reset(reset), .m_out(m_out2), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out2), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod3(.clk(clk), .reset(reset), .m_out(m_out3), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out3), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod4(.clk(clk), .reset(reset), .m_out(m_out4), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out4), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod5(.clk(clk), .reset(reset), .m_out(m_out5), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out5), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod6(.clk(clk), .reset(reset), .m_out(m_out6), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out6), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	datapath #(16, 1) datapathMod7(.clk(clk), .reset(reset), .m_out(m_out7), .v_out(v_out),.en_acc(en_acc),
									.output_data(parallel_out7), .clear_acc(clear_acc), .output_valid(output_valid),
									.output_ready(output_ready));

	l3_fc3_16_12_16_1_8_W_rom  matrixRom(.clk(clk),.addr0(addr_w0), .addr1(addr_w1), .addr2(addr_w2), .addr3(addr_w3), .addr4(addr_w4), .addr5(addr_w5), .addr6(addr_w6), .addr7(addr_w7), .z0(m_out0), .z1(m_out1), .z2(m_out2), .z3(m_out3), .z4(m_out4), .z5(m_out5), .z6(m_out6), .z7(m_out7));

endmodule

module l3_fc3_16_12_16_1_8_mux(parallel_out0, parallel_out1, parallel_out2, parallel_out3, parallel_out4, parallel_out5, parallel_out6, parallel_out7, sel, f);
	parameter T = 16;
	parameter P = 8;

	output signed [T-1 : 0] f;
	input logic unsigned [2 : 0] sel;
	input signed [T-1 : 0] parallel_out0;
	input signed [T-1 : 0] parallel_out1;
	input signed [T-1 : 0] parallel_out2;
	input signed [T-1 : 0] parallel_out3;
	input signed [T-1 : 0] parallel_out4;
	input signed [T-1 : 0] parallel_out5;
	input signed [T-1 : 0] parallel_out6;
	input signed [T-1 : 0] parallel_out7;
	logic unsigned [P*T-1 : 0] array;
	assign  array = {parallel_out0[15 : 0], parallel_out1[15 : 0], parallel_out2[15 : 0], parallel_out3[15 : 0], parallel_out4[15 : 0], parallel_out5[15 : 0], parallel_out6[15 : 0], parallel_out7[15: 0]};

	assign f = (sel == 0) ? parallel_out0 : 
			(sel == 1) ? parallel_out1 : 
			(sel == 2) ? parallel_out2 : 
			(sel == 3) ? parallel_out3 : 
			(sel == 4) ? parallel_out4 : 
			(sel == 5) ? parallel_out5 : 
			(sel == 6) ? parallel_out6 : 
			(sel == 7) ? parallel_out7 : 16'b0;
endmodule

module l3_fc3_16_12_16_1_8_W_rom(clk, addr0, addr1, addr2, addr3, addr4, addr5, addr6, addr7, z0, z1, z2, z3, z4, z5, z6, z7);
	input clk;
	input [7:0] addr0;
	input [7:0] addr1;
	input [7:0] addr2;
	input [7:0] addr3;
	input [7:0] addr4;
	input [7:0] addr5;
	input [7:0] addr6;
	input [7:0] addr7;
	output logic signed [15:0] z0;
	output logic signed [15:0] z1;
	output logic signed [15:0] z2;
	output logic signed [15:0] z3;
	output logic signed [15:0] z4;
	output logic signed [15:0] z5;
	output logic signed [15:0] z6;
	output logic signed [15:0] z7;
	always_ff @(posedge clk) begin
		case(addr0)
		0: z0 <= 16'd7;
		1: z0 <= 16'd5;
		2: z0 <= 16'd0;
		3: z0 <= -16'd5;
		4: z0 <= 16'd1;
		5: z0 <= 16'd7;
		6: z0 <= 16'd4;
		7: z0 <= 16'd0;
		8: z0 <= 16'd7;
		9: z0 <= -16'd3;
		10: z0 <= 16'd5;
		11: z0 <= -16'd5;
		12: z0 <= 16'd2;
		13: z0 <= -16'd3;
		14: z0 <= -16'd6;
		15: z0 <= -16'd7;
		16: z0 <= -16'd8;
		17: z0 <= -16'd3;
		18: z0 <= -16'd2;
		19: z0 <= -16'd4;
		20: z0 <= 16'd0;
		21: z0 <= 16'd1;
		22: z0 <= -16'd7;
		23: z0 <= -16'd8;
		24: z0 <= 16'd6;
		25: z0 <= 16'd0;
		26: z0 <= -16'd2;
		27: z0 <= 16'd0;
		28: z0 <= -16'd6;
		29: z0 <= -16'd6;
		30: z0 <= 16'd4;
		31: z0 <= -16'd7;
		32: z0 <= 16'd7;
		33: z0 <= -16'd4;
		34: z0 <= -16'd4;
		35: z0 <= 16'd1;
		36: z0 <= -16'd4;
		37: z0 <= -16'd8;
		38: z0 <= -16'd7;
		39: z0 <= -16'd5;
		40: z0 <= -16'd2;
		41: z0 <= 16'd6;
		42: z0 <= -16'd2;
		43: z0 <= -16'd8;
		44: z0 <= -16'd4;
		45: z0 <= 16'd0;
		46: z0 <= -16'd7;
		47: z0 <= -16'd4;
		48: z0 <= 16'd5;
		49: z0 <= -16'd1;
		50: z0 <= 16'd0;
		51: z0 <= -16'd2;
		52: z0 <= -16'd7;
		53: z0 <= 16'd1;
		54: z0 <= -16'd2;
		55: z0 <= 16'd7;
		56: z0 <= -16'd7;
		57: z0 <= 16'd4;
		58: z0 <= -16'd1;
		59: z0 <= -16'd5;
		60: z0 <= 16'd6;
		61: z0 <= -16'd5;
		62: z0 <= -16'd4;
		63: z0 <= 16'd5;
		64: z0 <= 16'd0;
		65: z0 <= 16'd1;
		66: z0 <= -16'd2;
		67: z0 <= 16'd4;
		68: z0 <= 16'd1;
		69: z0 <= 16'd0;
		70: z0 <= 16'd7;
		71: z0 <= 16'd7;
		72: z0 <= -16'd2;
		73: z0 <= -16'd3;
		74: z0 <= -16'd8;
		75: z0 <= 16'd2;
		76: z0 <= 16'd5;
		77: z0 <= -16'd7;
		78: z0 <= 16'd6;
		79: z0 <= 16'd2;
		80: z0 <= 16'd1;
		81: z0 <= -16'd1;
		82: z0 <= -16'd8;
		83: z0 <= 16'd2;
		84: z0 <= -16'd8;
		85: z0 <= -16'd2;
		86: z0 <= 16'd1;
		87: z0 <= -16'd6;
		88: z0 <= -16'd6;
		89: z0 <= -16'd7;
		90: z0 <= -16'd3;
		91: z0 <= -16'd8;
		92: z0 <= -16'd4;
		93: z0 <= 16'd2;
		94: z0 <= 16'd6;
		95: z0 <= 16'd4;
		96: z0 <= -16'd5;
		97: z0 <= -16'd4;
		98: z0 <= 16'd0;
		99: z0 <= 16'd4;
		100: z0 <= 16'd4;
		101: z0 <= -16'd1;
		102: z0 <= 16'd4;
		103: z0 <= -16'd5;
		104: z0 <= 16'd4;
		105: z0 <= 16'd4;
		106: z0 <= 16'd5;
		107: z0 <= 16'd1;
		108: z0 <= 16'd5;
		109: z0 <= 16'd4;
		110: z0 <= -16'd4;
		111: z0 <= -16'd2;
		112: z0 <= -16'd5;
		113: z0 <= -16'd4;
		114: z0 <= -16'd8;
		115: z0 <= -16'd5;
		116: z0 <= 16'd3;
		117: z0 <= 16'd2;
		118: z0 <= -16'd3;
		119: z0 <= 16'd5;
		120: z0 <= 16'd3;
		121: z0 <= 16'd3;
		122: z0 <= 16'd6;
		123: z0 <= 16'd7;
		124: z0 <= -16'd3;
		125: z0 <= 16'd4;
		126: z0 <= 16'd4;
		127: z0 <= 16'd0;
		128: z0 <= -16'd8;
		129: z0 <= -16'd4;
		130: z0 <= -16'd4;
		131: z0 <= 16'd5;
		132: z0 <= 16'd4;
		133: z0 <= -16'd8;
		134: z0 <= -16'd8;
		135: z0 <= 16'd0;
		136: z0 <= 16'd4;
		137: z0 <= 16'd5;
		138: z0 <= -16'd6;
		139: z0 <= 16'd2;
		140: z0 <= 16'd1;
		141: z0 <= -16'd2;
		142: z0 <= -16'd8;
		143: z0 <= 16'd4;
		144: z0 <= 16'd2;
		145: z0 <= -16'd7;
		146: z0 <= -16'd8;
		147: z0 <= -16'd3;
		148: z0 <= 16'd3;
		149: z0 <= -16'd3;
		150: z0 <= -16'd5;
		151: z0 <= -16'd2;
		152: z0 <= -16'd8;
		153: z0 <= -16'd7;
		154: z0 <= -16'd3;
		155: z0 <= -16'd3;
		156: z0 <= 16'd5;
		157: z0 <= -16'd7;
		158: z0 <= 16'd5;
		159: z0 <= 16'd5;
		160: z0 <= -16'd2;
		161: z0 <= -16'd6;
		162: z0 <= 16'd2;
		163: z0 <= -16'd6;
		164: z0 <= -16'd6;
		165: z0 <= 16'd2;
		166: z0 <= 16'd2;
		167: z0 <= 16'd7;
		168: z0 <= 16'd0;
		169: z0 <= 16'd4;
		170: z0 <= 16'd1;
		171: z0 <= -16'd7;
		172: z0 <= -16'd6;
		173: z0 <= 16'd1;
		174: z0 <= 16'd6;
		175: z0 <= 16'd5;
		176: z0 <= 16'd2;
		177: z0 <= 16'd6;
		178: z0 <= -16'd6;
		179: z0 <= -16'd3;
		180: z0 <= -16'd5;
		181: z0 <= -16'd3;
		182: z0 <= 16'd3;
		183: z0 <= -16'd4;
		184: z0 <= -16'd2;
		185: z0 <= -16'd7;
		186: z0 <= 16'd1;
		187: z0 <= -16'd5;
		188: z0 <= -16'd6;
		189: z0 <= -16'd1;
		190: z0 <= -16'd7;
		191: z0 <= 16'd0;
		endcase
		case(addr1)
		0: z1 <= 16'd7;
		1: z1 <= 16'd5;
		2: z1 <= 16'd0;
		3: z1 <= -16'd5;
		4: z1 <= 16'd1;
		5: z1 <= 16'd7;
		6: z1 <= 16'd4;
		7: z1 <= 16'd0;
		8: z1 <= 16'd7;
		9: z1 <= -16'd3;
		10: z1 <= 16'd5;
		11: z1 <= -16'd5;
		12: z1 <= 16'd2;
		13: z1 <= -16'd3;
		14: z1 <= -16'd6;
		15: z1 <= -16'd7;
		16: z1 <= -16'd8;
		17: z1 <= -16'd3;
		18: z1 <= -16'd2;
		19: z1 <= -16'd4;
		20: z1 <= 16'd0;
		21: z1 <= 16'd1;
		22: z1 <= -16'd7;
		23: z1 <= -16'd8;
		24: z1 <= 16'd6;
		25: z1 <= 16'd0;
		26: z1 <= -16'd2;
		27: z1 <= 16'd0;
		28: z1 <= -16'd6;
		29: z1 <= -16'd6;
		30: z1 <= 16'd4;
		31: z1 <= -16'd7;
		32: z1 <= 16'd7;
		33: z1 <= -16'd4;
		34: z1 <= -16'd4;
		35: z1 <= 16'd1;
		36: z1 <= -16'd4;
		37: z1 <= -16'd8;
		38: z1 <= -16'd7;
		39: z1 <= -16'd5;
		40: z1 <= -16'd2;
		41: z1 <= 16'd6;
		42: z1 <= -16'd2;
		43: z1 <= -16'd8;
		44: z1 <= -16'd4;
		45: z1 <= 16'd0;
		46: z1 <= -16'd7;
		47: z1 <= -16'd4;
		48: z1 <= 16'd5;
		49: z1 <= -16'd1;
		50: z1 <= 16'd0;
		51: z1 <= -16'd2;
		52: z1 <= -16'd7;
		53: z1 <= 16'd1;
		54: z1 <= -16'd2;
		55: z1 <= 16'd7;
		56: z1 <= -16'd7;
		57: z1 <= 16'd4;
		58: z1 <= -16'd1;
		59: z1 <= -16'd5;
		60: z1 <= 16'd6;
		61: z1 <= -16'd5;
		62: z1 <= -16'd4;
		63: z1 <= 16'd5;
		64: z1 <= 16'd0;
		65: z1 <= 16'd1;
		66: z1 <= -16'd2;
		67: z1 <= 16'd4;
		68: z1 <= 16'd1;
		69: z1 <= 16'd0;
		70: z1 <= 16'd7;
		71: z1 <= 16'd7;
		72: z1 <= -16'd2;
		73: z1 <= -16'd3;
		74: z1 <= -16'd8;
		75: z1 <= 16'd2;
		76: z1 <= 16'd5;
		77: z1 <= -16'd7;
		78: z1 <= 16'd6;
		79: z1 <= 16'd2;
		80: z1 <= 16'd1;
		81: z1 <= -16'd1;
		82: z1 <= -16'd8;
		83: z1 <= 16'd2;
		84: z1 <= -16'd8;
		85: z1 <= -16'd2;
		86: z1 <= 16'd1;
		87: z1 <= -16'd6;
		88: z1 <= -16'd6;
		89: z1 <= -16'd7;
		90: z1 <= -16'd3;
		91: z1 <= -16'd8;
		92: z1 <= -16'd4;
		93: z1 <= 16'd2;
		94: z1 <= 16'd6;
		95: z1 <= 16'd4;
		96: z1 <= -16'd5;
		97: z1 <= -16'd4;
		98: z1 <= 16'd0;
		99: z1 <= 16'd4;
		100: z1 <= 16'd4;
		101: z1 <= -16'd1;
		102: z1 <= 16'd4;
		103: z1 <= -16'd5;
		104: z1 <= 16'd4;
		105: z1 <= 16'd4;
		106: z1 <= 16'd5;
		107: z1 <= 16'd1;
		108: z1 <= 16'd5;
		109: z1 <= 16'd4;
		110: z1 <= -16'd4;
		111: z1 <= -16'd2;
		112: z1 <= -16'd5;
		113: z1 <= -16'd4;
		114: z1 <= -16'd8;
		115: z1 <= -16'd5;
		116: z1 <= 16'd3;
		117: z1 <= 16'd2;
		118: z1 <= -16'd3;
		119: z1 <= 16'd5;
		120: z1 <= 16'd3;
		121: z1 <= 16'd3;
		122: z1 <= 16'd6;
		123: z1 <= 16'd7;
		124: z1 <= -16'd3;
		125: z1 <= 16'd4;
		126: z1 <= 16'd4;
		127: z1 <= 16'd0;
		128: z1 <= -16'd8;
		129: z1 <= -16'd4;
		130: z1 <= -16'd4;
		131: z1 <= 16'd5;
		132: z1 <= 16'd4;
		133: z1 <= -16'd8;
		134: z1 <= -16'd8;
		135: z1 <= 16'd0;
		136: z1 <= 16'd4;
		137: z1 <= 16'd5;
		138: z1 <= -16'd6;
		139: z1 <= 16'd2;
		140: z1 <= 16'd1;
		141: z1 <= -16'd2;
		142: z1 <= -16'd8;
		143: z1 <= 16'd4;
		144: z1 <= 16'd2;
		145: z1 <= -16'd7;
		146: z1 <= -16'd8;
		147: z1 <= -16'd3;
		148: z1 <= 16'd3;
		149: z1 <= -16'd3;
		150: z1 <= -16'd5;
		151: z1 <= -16'd2;
		152: z1 <= -16'd8;
		153: z1 <= -16'd7;
		154: z1 <= -16'd3;
		155: z1 <= -16'd3;
		156: z1 <= 16'd5;
		157: z1 <= -16'd7;
		158: z1 <= 16'd5;
		159: z1 <= 16'd5;
		160: z1 <= -16'd2;
		161: z1 <= -16'd6;
		162: z1 <= 16'd2;
		163: z1 <= -16'd6;
		164: z1 <= -16'd6;
		165: z1 <= 16'd2;
		166: z1 <= 16'd2;
		167: z1 <= 16'd7;
		168: z1 <= 16'd0;
		169: z1 <= 16'd4;
		170: z1 <= 16'd1;
		171: z1 <= -16'd7;
		172: z1 <= -16'd6;
		173: z1 <= 16'd1;
		174: z1 <= 16'd6;
		175: z1 <= 16'd5;
		176: z1 <= 16'd2;
		177: z1 <= 16'd6;
		178: z1 <= -16'd6;
		179: z1 <= -16'd3;
		180: z1 <= -16'd5;
		181: z1 <= -16'd3;
		182: z1 <= 16'd3;
		183: z1 <= -16'd4;
		184: z1 <= -16'd2;
		185: z1 <= -16'd7;
		186: z1 <= 16'd1;
		187: z1 <= -16'd5;
		188: z1 <= -16'd6;
		189: z1 <= -16'd1;
		190: z1 <= -16'd7;
		191: z1 <= 16'd0;
		endcase
		case(addr2)
		0: z2 <= 16'd7;
		1: z2 <= 16'd5;
		2: z2 <= 16'd0;
		3: z2 <= -16'd5;
		4: z2 <= 16'd1;
		5: z2 <= 16'd7;
		6: z2 <= 16'd4;
		7: z2 <= 16'd0;
		8: z2 <= 16'd7;
		9: z2 <= -16'd3;
		10: z2 <= 16'd5;
		11: z2 <= -16'd5;
		12: z2 <= 16'd2;
		13: z2 <= -16'd3;
		14: z2 <= -16'd6;
		15: z2 <= -16'd7;
		16: z2 <= -16'd8;
		17: z2 <= -16'd3;
		18: z2 <= -16'd2;
		19: z2 <= -16'd4;
		20: z2 <= 16'd0;
		21: z2 <= 16'd1;
		22: z2 <= -16'd7;
		23: z2 <= -16'd8;
		24: z2 <= 16'd6;
		25: z2 <= 16'd0;
		26: z2 <= -16'd2;
		27: z2 <= 16'd0;
		28: z2 <= -16'd6;
		29: z2 <= -16'd6;
		30: z2 <= 16'd4;
		31: z2 <= -16'd7;
		32: z2 <= 16'd7;
		33: z2 <= -16'd4;
		34: z2 <= -16'd4;
		35: z2 <= 16'd1;
		36: z2 <= -16'd4;
		37: z2 <= -16'd8;
		38: z2 <= -16'd7;
		39: z2 <= -16'd5;
		40: z2 <= -16'd2;
		41: z2 <= 16'd6;
		42: z2 <= -16'd2;
		43: z2 <= -16'd8;
		44: z2 <= -16'd4;
		45: z2 <= 16'd0;
		46: z2 <= -16'd7;
		47: z2 <= -16'd4;
		48: z2 <= 16'd5;
		49: z2 <= -16'd1;
		50: z2 <= 16'd0;
		51: z2 <= -16'd2;
		52: z2 <= -16'd7;
		53: z2 <= 16'd1;
		54: z2 <= -16'd2;
		55: z2 <= 16'd7;
		56: z2 <= -16'd7;
		57: z2 <= 16'd4;
		58: z2 <= -16'd1;
		59: z2 <= -16'd5;
		60: z2 <= 16'd6;
		61: z2 <= -16'd5;
		62: z2 <= -16'd4;
		63: z2 <= 16'd5;
		64: z2 <= 16'd0;
		65: z2 <= 16'd1;
		66: z2 <= -16'd2;
		67: z2 <= 16'd4;
		68: z2 <= 16'd1;
		69: z2 <= 16'd0;
		70: z2 <= 16'd7;
		71: z2 <= 16'd7;
		72: z2 <= -16'd2;
		73: z2 <= -16'd3;
		74: z2 <= -16'd8;
		75: z2 <= 16'd2;
		76: z2 <= 16'd5;
		77: z2 <= -16'd7;
		78: z2 <= 16'd6;
		79: z2 <= 16'd2;
		80: z2 <= 16'd1;
		81: z2 <= -16'd1;
		82: z2 <= -16'd8;
		83: z2 <= 16'd2;
		84: z2 <= -16'd8;
		85: z2 <= -16'd2;
		86: z2 <= 16'd1;
		87: z2 <= -16'd6;
		88: z2 <= -16'd6;
		89: z2 <= -16'd7;
		90: z2 <= -16'd3;
		91: z2 <= -16'd8;
		92: z2 <= -16'd4;
		93: z2 <= 16'd2;
		94: z2 <= 16'd6;
		95: z2 <= 16'd4;
		96: z2 <= -16'd5;
		97: z2 <= -16'd4;
		98: z2 <= 16'd0;
		99: z2 <= 16'd4;
		100: z2 <= 16'd4;
		101: z2 <= -16'd1;
		102: z2 <= 16'd4;
		103: z2 <= -16'd5;
		104: z2 <= 16'd4;
		105: z2 <= 16'd4;
		106: z2 <= 16'd5;
		107: z2 <= 16'd1;
		108: z2 <= 16'd5;
		109: z2 <= 16'd4;
		110: z2 <= -16'd4;
		111: z2 <= -16'd2;
		112: z2 <= -16'd5;
		113: z2 <= -16'd4;
		114: z2 <= -16'd8;
		115: z2 <= -16'd5;
		116: z2 <= 16'd3;
		117: z2 <= 16'd2;
		118: z2 <= -16'd3;
		119: z2 <= 16'd5;
		120: z2 <= 16'd3;
		121: z2 <= 16'd3;
		122: z2 <= 16'd6;
		123: z2 <= 16'd7;
		124: z2 <= -16'd3;
		125: z2 <= 16'd4;
		126: z2 <= 16'd4;
		127: z2 <= 16'd0;
		128: z2 <= -16'd8;
		129: z2 <= -16'd4;
		130: z2 <= -16'd4;
		131: z2 <= 16'd5;
		132: z2 <= 16'd4;
		133: z2 <= -16'd8;
		134: z2 <= -16'd8;
		135: z2 <= 16'd0;
		136: z2 <= 16'd4;
		137: z2 <= 16'd5;
		138: z2 <= -16'd6;
		139: z2 <= 16'd2;
		140: z2 <= 16'd1;
		141: z2 <= -16'd2;
		142: z2 <= -16'd8;
		143: z2 <= 16'd4;
		144: z2 <= 16'd2;
		145: z2 <= -16'd7;
		146: z2 <= -16'd8;
		147: z2 <= -16'd3;
		148: z2 <= 16'd3;
		149: z2 <= -16'd3;
		150: z2 <= -16'd5;
		151: z2 <= -16'd2;
		152: z2 <= -16'd8;
		153: z2 <= -16'd7;
		154: z2 <= -16'd3;
		155: z2 <= -16'd3;
		156: z2 <= 16'd5;
		157: z2 <= -16'd7;
		158: z2 <= 16'd5;
		159: z2 <= 16'd5;
		160: z2 <= -16'd2;
		161: z2 <= -16'd6;
		162: z2 <= 16'd2;
		163: z2 <= -16'd6;
		164: z2 <= -16'd6;
		165: z2 <= 16'd2;
		166: z2 <= 16'd2;
		167: z2 <= 16'd7;
		168: z2 <= 16'd0;
		169: z2 <= 16'd4;
		170: z2 <= 16'd1;
		171: z2 <= -16'd7;
		172: z2 <= -16'd6;
		173: z2 <= 16'd1;
		174: z2 <= 16'd6;
		175: z2 <= 16'd5;
		176: z2 <= 16'd2;
		177: z2 <= 16'd6;
		178: z2 <= -16'd6;
		179: z2 <= -16'd3;
		180: z2 <= -16'd5;
		181: z2 <= -16'd3;
		182: z2 <= 16'd3;
		183: z2 <= -16'd4;
		184: z2 <= -16'd2;
		185: z2 <= -16'd7;
		186: z2 <= 16'd1;
		187: z2 <= -16'd5;
		188: z2 <= -16'd6;
		189: z2 <= -16'd1;
		190: z2 <= -16'd7;
		191: z2 <= 16'd0;
		endcase
		case(addr3)
		0: z3 <= 16'd7;
		1: z3 <= 16'd5;
		2: z3 <= 16'd0;
		3: z3 <= -16'd5;
		4: z3 <= 16'd1;
		5: z3 <= 16'd7;
		6: z3 <= 16'd4;
		7: z3 <= 16'd0;
		8: z3 <= 16'd7;
		9: z3 <= -16'd3;
		10: z3 <= 16'd5;
		11: z3 <= -16'd5;
		12: z3 <= 16'd2;
		13: z3 <= -16'd3;
		14: z3 <= -16'd6;
		15: z3 <= -16'd7;
		16: z3 <= -16'd8;
		17: z3 <= -16'd3;
		18: z3 <= -16'd2;
		19: z3 <= -16'd4;
		20: z3 <= 16'd0;
		21: z3 <= 16'd1;
		22: z3 <= -16'd7;
		23: z3 <= -16'd8;
		24: z3 <= 16'd6;
		25: z3 <= 16'd0;
		26: z3 <= -16'd2;
		27: z3 <= 16'd0;
		28: z3 <= -16'd6;
		29: z3 <= -16'd6;
		30: z3 <= 16'd4;
		31: z3 <= -16'd7;
		32: z3 <= 16'd7;
		33: z3 <= -16'd4;
		34: z3 <= -16'd4;
		35: z3 <= 16'd1;
		36: z3 <= -16'd4;
		37: z3 <= -16'd8;
		38: z3 <= -16'd7;
		39: z3 <= -16'd5;
		40: z3 <= -16'd2;
		41: z3 <= 16'd6;
		42: z3 <= -16'd2;
		43: z3 <= -16'd8;
		44: z3 <= -16'd4;
		45: z3 <= 16'd0;
		46: z3 <= -16'd7;
		47: z3 <= -16'd4;
		48: z3 <= 16'd5;
		49: z3 <= -16'd1;
		50: z3 <= 16'd0;
		51: z3 <= -16'd2;
		52: z3 <= -16'd7;
		53: z3 <= 16'd1;
		54: z3 <= -16'd2;
		55: z3 <= 16'd7;
		56: z3 <= -16'd7;
		57: z3 <= 16'd4;
		58: z3 <= -16'd1;
		59: z3 <= -16'd5;
		60: z3 <= 16'd6;
		61: z3 <= -16'd5;
		62: z3 <= -16'd4;
		63: z3 <= 16'd5;
		64: z3 <= 16'd0;
		65: z3 <= 16'd1;
		66: z3 <= -16'd2;
		67: z3 <= 16'd4;
		68: z3 <= 16'd1;
		69: z3 <= 16'd0;
		70: z3 <= 16'd7;
		71: z3 <= 16'd7;
		72: z3 <= -16'd2;
		73: z3 <= -16'd3;
		74: z3 <= -16'd8;
		75: z3 <= 16'd2;
		76: z3 <= 16'd5;
		77: z3 <= -16'd7;
		78: z3 <= 16'd6;
		79: z3 <= 16'd2;
		80: z3 <= 16'd1;
		81: z3 <= -16'd1;
		82: z3 <= -16'd8;
		83: z3 <= 16'd2;
		84: z3 <= -16'd8;
		85: z3 <= -16'd2;
		86: z3 <= 16'd1;
		87: z3 <= -16'd6;
		88: z3 <= -16'd6;
		89: z3 <= -16'd7;
		90: z3 <= -16'd3;
		91: z3 <= -16'd8;
		92: z3 <= -16'd4;
		93: z3 <= 16'd2;
		94: z3 <= 16'd6;
		95: z3 <= 16'd4;
		96: z3 <= -16'd5;
		97: z3 <= -16'd4;
		98: z3 <= 16'd0;
		99: z3 <= 16'd4;
		100: z3 <= 16'd4;
		101: z3 <= -16'd1;
		102: z3 <= 16'd4;
		103: z3 <= -16'd5;
		104: z3 <= 16'd4;
		105: z3 <= 16'd4;
		106: z3 <= 16'd5;
		107: z3 <= 16'd1;
		108: z3 <= 16'd5;
		109: z3 <= 16'd4;
		110: z3 <= -16'd4;
		111: z3 <= -16'd2;
		112: z3 <= -16'd5;
		113: z3 <= -16'd4;
		114: z3 <= -16'd8;
		115: z3 <= -16'd5;
		116: z3 <= 16'd3;
		117: z3 <= 16'd2;
		118: z3 <= -16'd3;
		119: z3 <= 16'd5;
		120: z3 <= 16'd3;
		121: z3 <= 16'd3;
		122: z3 <= 16'd6;
		123: z3 <= 16'd7;
		124: z3 <= -16'd3;
		125: z3 <= 16'd4;
		126: z3 <= 16'd4;
		127: z3 <= 16'd0;
		128: z3 <= -16'd8;
		129: z3 <= -16'd4;
		130: z3 <= -16'd4;
		131: z3 <= 16'd5;
		132: z3 <= 16'd4;
		133: z3 <= -16'd8;
		134: z3 <= -16'd8;
		135: z3 <= 16'd0;
		136: z3 <= 16'd4;
		137: z3 <= 16'd5;
		138: z3 <= -16'd6;
		139: z3 <= 16'd2;
		140: z3 <= 16'd1;
		141: z3 <= -16'd2;
		142: z3 <= -16'd8;
		143: z3 <= 16'd4;
		144: z3 <= 16'd2;
		145: z3 <= -16'd7;
		146: z3 <= -16'd8;
		147: z3 <= -16'd3;
		148: z3 <= 16'd3;
		149: z3 <= -16'd3;
		150: z3 <= -16'd5;
		151: z3 <= -16'd2;
		152: z3 <= -16'd8;
		153: z3 <= -16'd7;
		154: z3 <= -16'd3;
		155: z3 <= -16'd3;
		156: z3 <= 16'd5;
		157: z3 <= -16'd7;
		158: z3 <= 16'd5;
		159: z3 <= 16'd5;
		160: z3 <= -16'd2;
		161: z3 <= -16'd6;
		162: z3 <= 16'd2;
		163: z3 <= -16'd6;
		164: z3 <= -16'd6;
		165: z3 <= 16'd2;
		166: z3 <= 16'd2;
		167: z3 <= 16'd7;
		168: z3 <= 16'd0;
		169: z3 <= 16'd4;
		170: z3 <= 16'd1;
		171: z3 <= -16'd7;
		172: z3 <= -16'd6;
		173: z3 <= 16'd1;
		174: z3 <= 16'd6;
		175: z3 <= 16'd5;
		176: z3 <= 16'd2;
		177: z3 <= 16'd6;
		178: z3 <= -16'd6;
		179: z3 <= -16'd3;
		180: z3 <= -16'd5;
		181: z3 <= -16'd3;
		182: z3 <= 16'd3;
		183: z3 <= -16'd4;
		184: z3 <= -16'd2;
		185: z3 <= -16'd7;
		186: z3 <= 16'd1;
		187: z3 <= -16'd5;
		188: z3 <= -16'd6;
		189: z3 <= -16'd1;
		190: z3 <= -16'd7;
		191: z3 <= 16'd0;
		endcase
		case(addr4)
		0: z4 <= 16'd7;
		1: z4 <= 16'd5;
		2: z4 <= 16'd0;
		3: z4 <= -16'd5;
		4: z4 <= 16'd1;
		5: z4 <= 16'd7;
		6: z4 <= 16'd4;
		7: z4 <= 16'd0;
		8: z4 <= 16'd7;
		9: z4 <= -16'd3;
		10: z4 <= 16'd5;
		11: z4 <= -16'd5;
		12: z4 <= 16'd2;
		13: z4 <= -16'd3;
		14: z4 <= -16'd6;
		15: z4 <= -16'd7;
		16: z4 <= -16'd8;
		17: z4 <= -16'd3;
		18: z4 <= -16'd2;
		19: z4 <= -16'd4;
		20: z4 <= 16'd0;
		21: z4 <= 16'd1;
		22: z4 <= -16'd7;
		23: z4 <= -16'd8;
		24: z4 <= 16'd6;
		25: z4 <= 16'd0;
		26: z4 <= -16'd2;
		27: z4 <= 16'd0;
		28: z4 <= -16'd6;
		29: z4 <= -16'd6;
		30: z4 <= 16'd4;
		31: z4 <= -16'd7;
		32: z4 <= 16'd7;
		33: z4 <= -16'd4;
		34: z4 <= -16'd4;
		35: z4 <= 16'd1;
		36: z4 <= -16'd4;
		37: z4 <= -16'd8;
		38: z4 <= -16'd7;
		39: z4 <= -16'd5;
		40: z4 <= -16'd2;
		41: z4 <= 16'd6;
		42: z4 <= -16'd2;
		43: z4 <= -16'd8;
		44: z4 <= -16'd4;
		45: z4 <= 16'd0;
		46: z4 <= -16'd7;
		47: z4 <= -16'd4;
		48: z4 <= 16'd5;
		49: z4 <= -16'd1;
		50: z4 <= 16'd0;
		51: z4 <= -16'd2;
		52: z4 <= -16'd7;
		53: z4 <= 16'd1;
		54: z4 <= -16'd2;
		55: z4 <= 16'd7;
		56: z4 <= -16'd7;
		57: z4 <= 16'd4;
		58: z4 <= -16'd1;
		59: z4 <= -16'd5;
		60: z4 <= 16'd6;
		61: z4 <= -16'd5;
		62: z4 <= -16'd4;
		63: z4 <= 16'd5;
		64: z4 <= 16'd0;
		65: z4 <= 16'd1;
		66: z4 <= -16'd2;
		67: z4 <= 16'd4;
		68: z4 <= 16'd1;
		69: z4 <= 16'd0;
		70: z4 <= 16'd7;
		71: z4 <= 16'd7;
		72: z4 <= -16'd2;
		73: z4 <= -16'd3;
		74: z4 <= -16'd8;
		75: z4 <= 16'd2;
		76: z4 <= 16'd5;
		77: z4 <= -16'd7;
		78: z4 <= 16'd6;
		79: z4 <= 16'd2;
		80: z4 <= 16'd1;
		81: z4 <= -16'd1;
		82: z4 <= -16'd8;
		83: z4 <= 16'd2;
		84: z4 <= -16'd8;
		85: z4 <= -16'd2;
		86: z4 <= 16'd1;
		87: z4 <= -16'd6;
		88: z4 <= -16'd6;
		89: z4 <= -16'd7;
		90: z4 <= -16'd3;
		91: z4 <= -16'd8;
		92: z4 <= -16'd4;
		93: z4 <= 16'd2;
		94: z4 <= 16'd6;
		95: z4 <= 16'd4;
		96: z4 <= -16'd5;
		97: z4 <= -16'd4;
		98: z4 <= 16'd0;
		99: z4 <= 16'd4;
		100: z4 <= 16'd4;
		101: z4 <= -16'd1;
		102: z4 <= 16'd4;
		103: z4 <= -16'd5;
		104: z4 <= 16'd4;
		105: z4 <= 16'd4;
		106: z4 <= 16'd5;
		107: z4 <= 16'd1;
		108: z4 <= 16'd5;
		109: z4 <= 16'd4;
		110: z4 <= -16'd4;
		111: z4 <= -16'd2;
		112: z4 <= -16'd5;
		113: z4 <= -16'd4;
		114: z4 <= -16'd8;
		115: z4 <= -16'd5;
		116: z4 <= 16'd3;
		117: z4 <= 16'd2;
		118: z4 <= -16'd3;
		119: z4 <= 16'd5;
		120: z4 <= 16'd3;
		121: z4 <= 16'd3;
		122: z4 <= 16'd6;
		123: z4 <= 16'd7;
		124: z4 <= -16'd3;
		125: z4 <= 16'd4;
		126: z4 <= 16'd4;
		127: z4 <= 16'd0;
		128: z4 <= -16'd8;
		129: z4 <= -16'd4;
		130: z4 <= -16'd4;
		131: z4 <= 16'd5;
		132: z4 <= 16'd4;
		133: z4 <= -16'd8;
		134: z4 <= -16'd8;
		135: z4 <= 16'd0;
		136: z4 <= 16'd4;
		137: z4 <= 16'd5;
		138: z4 <= -16'd6;
		139: z4 <= 16'd2;
		140: z4 <= 16'd1;
		141: z4 <= -16'd2;
		142: z4 <= -16'd8;
		143: z4 <= 16'd4;
		144: z4 <= 16'd2;
		145: z4 <= -16'd7;
		146: z4 <= -16'd8;
		147: z4 <= -16'd3;
		148: z4 <= 16'd3;
		149: z4 <= -16'd3;
		150: z4 <= -16'd5;
		151: z4 <= -16'd2;
		152: z4 <= -16'd8;
		153: z4 <= -16'd7;
		154: z4 <= -16'd3;
		155: z4 <= -16'd3;
		156: z4 <= 16'd5;
		157: z4 <= -16'd7;
		158: z4 <= 16'd5;
		159: z4 <= 16'd5;
		160: z4 <= -16'd2;
		161: z4 <= -16'd6;
		162: z4 <= 16'd2;
		163: z4 <= -16'd6;
		164: z4 <= -16'd6;
		165: z4 <= 16'd2;
		166: z4 <= 16'd2;
		167: z4 <= 16'd7;
		168: z4 <= 16'd0;
		169: z4 <= 16'd4;
		170: z4 <= 16'd1;
		171: z4 <= -16'd7;
		172: z4 <= -16'd6;
		173: z4 <= 16'd1;
		174: z4 <= 16'd6;
		175: z4 <= 16'd5;
		176: z4 <= 16'd2;
		177: z4 <= 16'd6;
		178: z4 <= -16'd6;
		179: z4 <= -16'd3;
		180: z4 <= -16'd5;
		181: z4 <= -16'd3;
		182: z4 <= 16'd3;
		183: z4 <= -16'd4;
		184: z4 <= -16'd2;
		185: z4 <= -16'd7;
		186: z4 <= 16'd1;
		187: z4 <= -16'd5;
		188: z4 <= -16'd6;
		189: z4 <= -16'd1;
		190: z4 <= -16'd7;
		191: z4 <= 16'd0;
		endcase
		case(addr5)
		0: z5 <= 16'd7;
		1: z5 <= 16'd5;
		2: z5 <= 16'd0;
		3: z5 <= -16'd5;
		4: z5 <= 16'd1;
		5: z5 <= 16'd7;
		6: z5 <= 16'd4;
		7: z5 <= 16'd0;
		8: z5 <= 16'd7;
		9: z5 <= -16'd3;
		10: z5 <= 16'd5;
		11: z5 <= -16'd5;
		12: z5 <= 16'd2;
		13: z5 <= -16'd3;
		14: z5 <= -16'd6;
		15: z5 <= -16'd7;
		16: z5 <= -16'd8;
		17: z5 <= -16'd3;
		18: z5 <= -16'd2;
		19: z5 <= -16'd4;
		20: z5 <= 16'd0;
		21: z5 <= 16'd1;
		22: z5 <= -16'd7;
		23: z5 <= -16'd8;
		24: z5 <= 16'd6;
		25: z5 <= 16'd0;
		26: z5 <= -16'd2;
		27: z5 <= 16'd0;
		28: z5 <= -16'd6;
		29: z5 <= -16'd6;
		30: z5 <= 16'd4;
		31: z5 <= -16'd7;
		32: z5 <= 16'd7;
		33: z5 <= -16'd4;
		34: z5 <= -16'd4;
		35: z5 <= 16'd1;
		36: z5 <= -16'd4;
		37: z5 <= -16'd8;
		38: z5 <= -16'd7;
		39: z5 <= -16'd5;
		40: z5 <= -16'd2;
		41: z5 <= 16'd6;
		42: z5 <= -16'd2;
		43: z5 <= -16'd8;
		44: z5 <= -16'd4;
		45: z5 <= 16'd0;
		46: z5 <= -16'd7;
		47: z5 <= -16'd4;
		48: z5 <= 16'd5;
		49: z5 <= -16'd1;
		50: z5 <= 16'd0;
		51: z5 <= -16'd2;
		52: z5 <= -16'd7;
		53: z5 <= 16'd1;
		54: z5 <= -16'd2;
		55: z5 <= 16'd7;
		56: z5 <= -16'd7;
		57: z5 <= 16'd4;
		58: z5 <= -16'd1;
		59: z5 <= -16'd5;
		60: z5 <= 16'd6;
		61: z5 <= -16'd5;
		62: z5 <= -16'd4;
		63: z5 <= 16'd5;
		64: z5 <= 16'd0;
		65: z5 <= 16'd1;
		66: z5 <= -16'd2;
		67: z5 <= 16'd4;
		68: z5 <= 16'd1;
		69: z5 <= 16'd0;
		70: z5 <= 16'd7;
		71: z5 <= 16'd7;
		72: z5 <= -16'd2;
		73: z5 <= -16'd3;
		74: z5 <= -16'd8;
		75: z5 <= 16'd2;
		76: z5 <= 16'd5;
		77: z5 <= -16'd7;
		78: z5 <= 16'd6;
		79: z5 <= 16'd2;
		80: z5 <= 16'd1;
		81: z5 <= -16'd1;
		82: z5 <= -16'd8;
		83: z5 <= 16'd2;
		84: z5 <= -16'd8;
		85: z5 <= -16'd2;
		86: z5 <= 16'd1;
		87: z5 <= -16'd6;
		88: z5 <= -16'd6;
		89: z5 <= -16'd7;
		90: z5 <= -16'd3;
		91: z5 <= -16'd8;
		92: z5 <= -16'd4;
		93: z5 <= 16'd2;
		94: z5 <= 16'd6;
		95: z5 <= 16'd4;
		96: z5 <= -16'd5;
		97: z5 <= -16'd4;
		98: z5 <= 16'd0;
		99: z5 <= 16'd4;
		100: z5 <= 16'd4;
		101: z5 <= -16'd1;
		102: z5 <= 16'd4;
		103: z5 <= -16'd5;
		104: z5 <= 16'd4;
		105: z5 <= 16'd4;
		106: z5 <= 16'd5;
		107: z5 <= 16'd1;
		108: z5 <= 16'd5;
		109: z5 <= 16'd4;
		110: z5 <= -16'd4;
		111: z5 <= -16'd2;
		112: z5 <= -16'd5;
		113: z5 <= -16'd4;
		114: z5 <= -16'd8;
		115: z5 <= -16'd5;
		116: z5 <= 16'd3;
		117: z5 <= 16'd2;
		118: z5 <= -16'd3;
		119: z5 <= 16'd5;
		120: z5 <= 16'd3;
		121: z5 <= 16'd3;
		122: z5 <= 16'd6;
		123: z5 <= 16'd7;
		124: z5 <= -16'd3;
		125: z5 <= 16'd4;
		126: z5 <= 16'd4;
		127: z5 <= 16'd0;
		128: z5 <= -16'd8;
		129: z5 <= -16'd4;
		130: z5 <= -16'd4;
		131: z5 <= 16'd5;
		132: z5 <= 16'd4;
		133: z5 <= -16'd8;
		134: z5 <= -16'd8;
		135: z5 <= 16'd0;
		136: z5 <= 16'd4;
		137: z5 <= 16'd5;
		138: z5 <= -16'd6;
		139: z5 <= 16'd2;
		140: z5 <= 16'd1;
		141: z5 <= -16'd2;
		142: z5 <= -16'd8;
		143: z5 <= 16'd4;
		144: z5 <= 16'd2;
		145: z5 <= -16'd7;
		146: z5 <= -16'd8;
		147: z5 <= -16'd3;
		148: z5 <= 16'd3;
		149: z5 <= -16'd3;
		150: z5 <= -16'd5;
		151: z5 <= -16'd2;
		152: z5 <= -16'd8;
		153: z5 <= -16'd7;
		154: z5 <= -16'd3;
		155: z5 <= -16'd3;
		156: z5 <= 16'd5;
		157: z5 <= -16'd7;
		158: z5 <= 16'd5;
		159: z5 <= 16'd5;
		160: z5 <= -16'd2;
		161: z5 <= -16'd6;
		162: z5 <= 16'd2;
		163: z5 <= -16'd6;
		164: z5 <= -16'd6;
		165: z5 <= 16'd2;
		166: z5 <= 16'd2;
		167: z5 <= 16'd7;
		168: z5 <= 16'd0;
		169: z5 <= 16'd4;
		170: z5 <= 16'd1;
		171: z5 <= -16'd7;
		172: z5 <= -16'd6;
		173: z5 <= 16'd1;
		174: z5 <= 16'd6;
		175: z5 <= 16'd5;
		176: z5 <= 16'd2;
		177: z5 <= 16'd6;
		178: z5 <= -16'd6;
		179: z5 <= -16'd3;
		180: z5 <= -16'd5;
		181: z5 <= -16'd3;
		182: z5 <= 16'd3;
		183: z5 <= -16'd4;
		184: z5 <= -16'd2;
		185: z5 <= -16'd7;
		186: z5 <= 16'd1;
		187: z5 <= -16'd5;
		188: z5 <= -16'd6;
		189: z5 <= -16'd1;
		190: z5 <= -16'd7;
		191: z5 <= 16'd0;
		endcase
		case(addr6)
		0: z6 <= 16'd7;
		1: z6 <= 16'd5;
		2: z6 <= 16'd0;
		3: z6 <= -16'd5;
		4: z6 <= 16'd1;
		5: z6 <= 16'd7;
		6: z6 <= 16'd4;
		7: z6 <= 16'd0;
		8: z6 <= 16'd7;
		9: z6 <= -16'd3;
		10: z6 <= 16'd5;
		11: z6 <= -16'd5;
		12: z6 <= 16'd2;
		13: z6 <= -16'd3;
		14: z6 <= -16'd6;
		15: z6 <= -16'd7;
		16: z6 <= -16'd8;
		17: z6 <= -16'd3;
		18: z6 <= -16'd2;
		19: z6 <= -16'd4;
		20: z6 <= 16'd0;
		21: z6 <= 16'd1;
		22: z6 <= -16'd7;
		23: z6 <= -16'd8;
		24: z6 <= 16'd6;
		25: z6 <= 16'd0;
		26: z6 <= -16'd2;
		27: z6 <= 16'd0;
		28: z6 <= -16'd6;
		29: z6 <= -16'd6;
		30: z6 <= 16'd4;
		31: z6 <= -16'd7;
		32: z6 <= 16'd7;
		33: z6 <= -16'd4;
		34: z6 <= -16'd4;
		35: z6 <= 16'd1;
		36: z6 <= -16'd4;
		37: z6 <= -16'd8;
		38: z6 <= -16'd7;
		39: z6 <= -16'd5;
		40: z6 <= -16'd2;
		41: z6 <= 16'd6;
		42: z6 <= -16'd2;
		43: z6 <= -16'd8;
		44: z6 <= -16'd4;
		45: z6 <= 16'd0;
		46: z6 <= -16'd7;
		47: z6 <= -16'd4;
		48: z6 <= 16'd5;
		49: z6 <= -16'd1;
		50: z6 <= 16'd0;
		51: z6 <= -16'd2;
		52: z6 <= -16'd7;
		53: z6 <= 16'd1;
		54: z6 <= -16'd2;
		55: z6 <= 16'd7;
		56: z6 <= -16'd7;
		57: z6 <= 16'd4;
		58: z6 <= -16'd1;
		59: z6 <= -16'd5;
		60: z6 <= 16'd6;
		61: z6 <= -16'd5;
		62: z6 <= -16'd4;
		63: z6 <= 16'd5;
		64: z6 <= 16'd0;
		65: z6 <= 16'd1;
		66: z6 <= -16'd2;
		67: z6 <= 16'd4;
		68: z6 <= 16'd1;
		69: z6 <= 16'd0;
		70: z6 <= 16'd7;
		71: z6 <= 16'd7;
		72: z6 <= -16'd2;
		73: z6 <= -16'd3;
		74: z6 <= -16'd8;
		75: z6 <= 16'd2;
		76: z6 <= 16'd5;
		77: z6 <= -16'd7;
		78: z6 <= 16'd6;
		79: z6 <= 16'd2;
		80: z6 <= 16'd1;
		81: z6 <= -16'd1;
		82: z6 <= -16'd8;
		83: z6 <= 16'd2;
		84: z6 <= -16'd8;
		85: z6 <= -16'd2;
		86: z6 <= 16'd1;
		87: z6 <= -16'd6;
		88: z6 <= -16'd6;
		89: z6 <= -16'd7;
		90: z6 <= -16'd3;
		91: z6 <= -16'd8;
		92: z6 <= -16'd4;
		93: z6 <= 16'd2;
		94: z6 <= 16'd6;
		95: z6 <= 16'd4;
		96: z6 <= -16'd5;
		97: z6 <= -16'd4;
		98: z6 <= 16'd0;
		99: z6 <= 16'd4;
		100: z6 <= 16'd4;
		101: z6 <= -16'd1;
		102: z6 <= 16'd4;
		103: z6 <= -16'd5;
		104: z6 <= 16'd4;
		105: z6 <= 16'd4;
		106: z6 <= 16'd5;
		107: z6 <= 16'd1;
		108: z6 <= 16'd5;
		109: z6 <= 16'd4;
		110: z6 <= -16'd4;
		111: z6 <= -16'd2;
		112: z6 <= -16'd5;
		113: z6 <= -16'd4;
		114: z6 <= -16'd8;
		115: z6 <= -16'd5;
		116: z6 <= 16'd3;
		117: z6 <= 16'd2;
		118: z6 <= -16'd3;
		119: z6 <= 16'd5;
		120: z6 <= 16'd3;
		121: z6 <= 16'd3;
		122: z6 <= 16'd6;
		123: z6 <= 16'd7;
		124: z6 <= -16'd3;
		125: z6 <= 16'd4;
		126: z6 <= 16'd4;
		127: z6 <= 16'd0;
		128: z6 <= -16'd8;
		129: z6 <= -16'd4;
		130: z6 <= -16'd4;
		131: z6 <= 16'd5;
		132: z6 <= 16'd4;
		133: z6 <= -16'd8;
		134: z6 <= -16'd8;
		135: z6 <= 16'd0;
		136: z6 <= 16'd4;
		137: z6 <= 16'd5;
		138: z6 <= -16'd6;
		139: z6 <= 16'd2;
		140: z6 <= 16'd1;
		141: z6 <= -16'd2;
		142: z6 <= -16'd8;
		143: z6 <= 16'd4;
		144: z6 <= 16'd2;
		145: z6 <= -16'd7;
		146: z6 <= -16'd8;
		147: z6 <= -16'd3;
		148: z6 <= 16'd3;
		149: z6 <= -16'd3;
		150: z6 <= -16'd5;
		151: z6 <= -16'd2;
		152: z6 <= -16'd8;
		153: z6 <= -16'd7;
		154: z6 <= -16'd3;
		155: z6 <= -16'd3;
		156: z6 <= 16'd5;
		157: z6 <= -16'd7;
		158: z6 <= 16'd5;
		159: z6 <= 16'd5;
		160: z6 <= -16'd2;
		161: z6 <= -16'd6;
		162: z6 <= 16'd2;
		163: z6 <= -16'd6;
		164: z6 <= -16'd6;
		165: z6 <= 16'd2;
		166: z6 <= 16'd2;
		167: z6 <= 16'd7;
		168: z6 <= 16'd0;
		169: z6 <= 16'd4;
		170: z6 <= 16'd1;
		171: z6 <= -16'd7;
		172: z6 <= -16'd6;
		173: z6 <= 16'd1;
		174: z6 <= 16'd6;
		175: z6 <= 16'd5;
		176: z6 <= 16'd2;
		177: z6 <= 16'd6;
		178: z6 <= -16'd6;
		179: z6 <= -16'd3;
		180: z6 <= -16'd5;
		181: z6 <= -16'd3;
		182: z6 <= 16'd3;
		183: z6 <= -16'd4;
		184: z6 <= -16'd2;
		185: z6 <= -16'd7;
		186: z6 <= 16'd1;
		187: z6 <= -16'd5;
		188: z6 <= -16'd6;
		189: z6 <= -16'd1;
		190: z6 <= -16'd7;
		191: z6 <= 16'd0;
		endcase
		case(addr7)
		0: z7 <= 16'd7;
		1: z7 <= 16'd5;
		2: z7 <= 16'd0;
		3: z7 <= -16'd5;
		4: z7 <= 16'd1;
		5: z7 <= 16'd7;
		6: z7 <= 16'd4;
		7: z7 <= 16'd0;
		8: z7 <= 16'd7;
		9: z7 <= -16'd3;
		10: z7 <= 16'd5;
		11: z7 <= -16'd5;
		12: z7 <= 16'd2;
		13: z7 <= -16'd3;
		14: z7 <= -16'd6;
		15: z7 <= -16'd7;
		16: z7 <= -16'd8;
		17: z7 <= -16'd3;
		18: z7 <= -16'd2;
		19: z7 <= -16'd4;
		20: z7 <= 16'd0;
		21: z7 <= 16'd1;
		22: z7 <= -16'd7;
		23: z7 <= -16'd8;
		24: z7 <= 16'd6;
		25: z7 <= 16'd0;
		26: z7 <= -16'd2;
		27: z7 <= 16'd0;
		28: z7 <= -16'd6;
		29: z7 <= -16'd6;
		30: z7 <= 16'd4;
		31: z7 <= -16'd7;
		32: z7 <= 16'd7;
		33: z7 <= -16'd4;
		34: z7 <= -16'd4;
		35: z7 <= 16'd1;
		36: z7 <= -16'd4;
		37: z7 <= -16'd8;
		38: z7 <= -16'd7;
		39: z7 <= -16'd5;
		40: z7 <= -16'd2;
		41: z7 <= 16'd6;
		42: z7 <= -16'd2;
		43: z7 <= -16'd8;
		44: z7 <= -16'd4;
		45: z7 <= 16'd0;
		46: z7 <= -16'd7;
		47: z7 <= -16'd4;
		48: z7 <= 16'd5;
		49: z7 <= -16'd1;
		50: z7 <= 16'd0;
		51: z7 <= -16'd2;
		52: z7 <= -16'd7;
		53: z7 <= 16'd1;
		54: z7 <= -16'd2;
		55: z7 <= 16'd7;
		56: z7 <= -16'd7;
		57: z7 <= 16'd4;
		58: z7 <= -16'd1;
		59: z7 <= -16'd5;
		60: z7 <= 16'd6;
		61: z7 <= -16'd5;
		62: z7 <= -16'd4;
		63: z7 <= 16'd5;
		64: z7 <= 16'd0;
		65: z7 <= 16'd1;
		66: z7 <= -16'd2;
		67: z7 <= 16'd4;
		68: z7 <= 16'd1;
		69: z7 <= 16'd0;
		70: z7 <= 16'd7;
		71: z7 <= 16'd7;
		72: z7 <= -16'd2;
		73: z7 <= -16'd3;
		74: z7 <= -16'd8;
		75: z7 <= 16'd2;
		76: z7 <= 16'd5;
		77: z7 <= -16'd7;
		78: z7 <= 16'd6;
		79: z7 <= 16'd2;
		80: z7 <= 16'd1;
		81: z7 <= -16'd1;
		82: z7 <= -16'd8;
		83: z7 <= 16'd2;
		84: z7 <= -16'd8;
		85: z7 <= -16'd2;
		86: z7 <= 16'd1;
		87: z7 <= -16'd6;
		88: z7 <= -16'd6;
		89: z7 <= -16'd7;
		90: z7 <= -16'd3;
		91: z7 <= -16'd8;
		92: z7 <= -16'd4;
		93: z7 <= 16'd2;
		94: z7 <= 16'd6;
		95: z7 <= 16'd4;
		96: z7 <= -16'd5;
		97: z7 <= -16'd4;
		98: z7 <= 16'd0;
		99: z7 <= 16'd4;
		100: z7 <= 16'd4;
		101: z7 <= -16'd1;
		102: z7 <= 16'd4;
		103: z7 <= -16'd5;
		104: z7 <= 16'd4;
		105: z7 <= 16'd4;
		106: z7 <= 16'd5;
		107: z7 <= 16'd1;
		108: z7 <= 16'd5;
		109: z7 <= 16'd4;
		110: z7 <= -16'd4;
		111: z7 <= -16'd2;
		112: z7 <= -16'd5;
		113: z7 <= -16'd4;
		114: z7 <= -16'd8;
		115: z7 <= -16'd5;
		116: z7 <= 16'd3;
		117: z7 <= 16'd2;
		118: z7 <= -16'd3;
		119: z7 <= 16'd5;
		120: z7 <= 16'd3;
		121: z7 <= 16'd3;
		122: z7 <= 16'd6;
		123: z7 <= 16'd7;
		124: z7 <= -16'd3;
		125: z7 <= 16'd4;
		126: z7 <= 16'd4;
		127: z7 <= 16'd0;
		128: z7 <= -16'd8;
		129: z7 <= -16'd4;
		130: z7 <= -16'd4;
		131: z7 <= 16'd5;
		132: z7 <= 16'd4;
		133: z7 <= -16'd8;
		134: z7 <= -16'd8;
		135: z7 <= 16'd0;
		136: z7 <= 16'd4;
		137: z7 <= 16'd5;
		138: z7 <= -16'd6;
		139: z7 <= 16'd2;
		140: z7 <= 16'd1;
		141: z7 <= -16'd2;
		142: z7 <= -16'd8;
		143: z7 <= 16'd4;
		144: z7 <= 16'd2;
		145: z7 <= -16'd7;
		146: z7 <= -16'd8;
		147: z7 <= -16'd3;
		148: z7 <= 16'd3;
		149: z7 <= -16'd3;
		150: z7 <= -16'd5;
		151: z7 <= -16'd2;
		152: z7 <= -16'd8;
		153: z7 <= -16'd7;
		154: z7 <= -16'd3;
		155: z7 <= -16'd3;
		156: z7 <= 16'd5;
		157: z7 <= -16'd7;
		158: z7 <= 16'd5;
		159: z7 <= 16'd5;
		160: z7 <= -16'd2;
		161: z7 <= -16'd6;
		162: z7 <= 16'd2;
		163: z7 <= -16'd6;
		164: z7 <= -16'd6;
		165: z7 <= 16'd2;
		166: z7 <= 16'd2;
		167: z7 <= 16'd7;
		168: z7 <= 16'd0;
		169: z7 <= 16'd4;
		170: z7 <= 16'd1;
		171: z7 <= -16'd7;
		172: z7 <= -16'd6;
		173: z7 <= 16'd1;
		174: z7 <= 16'd6;
		175: z7 <= 16'd5;
		176: z7 <= 16'd2;
		177: z7 <= 16'd6;
		178: z7 <= -16'd6;
		179: z7 <= -16'd3;
		180: z7 <= -16'd5;
		181: z7 <= -16'd3;
		182: z7 <= 16'd3;
		183: z7 <= -16'd4;
		184: z7 <= -16'd2;
		185: z7 <= -16'd7;
		186: z7 <= 16'd1;
		187: z7 <= -16'd5;
		188: z7 <= -16'd6;
		189: z7 <= -16'd1;
		190: z7 <= -16'd7;
		191: z7 <= 16'd0;
		endcase
	end
endmodule

